memory_inst : memory PORT MAP (
		address	 => address_sig,
		data	 => data_sig,
		we	 => we_sig,
		q	 => q_sig
	);
