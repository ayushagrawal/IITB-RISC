library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;

package
