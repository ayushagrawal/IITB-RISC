// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 16.0.0 Build 211 04/27/2016 SJ Standard Edition"

// DATE "10/14/2016 22:55:27"

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module memory (
	address,
	data,
	we,
	q)/* synthesis synthesis_greybox=0 */;
input 	[4:0] address;
input 	[15:0] data;
input 	we;
output 	[15:0] q;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209_combout ;


memory_LPM_RAM_DQ_1 lpm_ram_dq_component(
	.address_0(address[0]),
	.address_1(address[1]),
	.address_2(address[2]),
	.address_4(address[4]),
	.address_3(address[3]),
	.result_node_0(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14_combout ),
	.result_node_1(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27_combout ),
	.result_node_2(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40_combout ),
	.result_node_3(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53_combout ),
	.result_node_4(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66_combout ),
	.result_node_5(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79_combout ),
	.result_node_6(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92_combout ),
	.result_node_7(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105_combout ),
	.result_node_8(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118_combout ),
	.result_node_9(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131_combout ),
	.result_node_10(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144_combout ),
	.result_node_11(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157_combout ),
	.result_node_12(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170_combout ),
	.result_node_13(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183_combout ),
	.result_node_14(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196_combout ),
	.result_node_15(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209_combout ),
	.data_0(data[0]),
	.we(we),
	.data_1(data[1]),
	.data_2(data[2]),
	.data_3(data[3]),
	.data_4(data[4]),
	.data_5(data[5]),
	.data_6(data[6]),
	.data_7(data[7]),
	.data_8(data[8]),
	.data_9(data[9]),
	.data_10(data[10]),
	.data_11(data[11]),
	.data_12(data[12]),
	.data_13(data[13]),
	.data_14(data[14]),
	.data_15(data[15]));

assign q[0] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14_combout ;

assign q[1] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27_combout ;

assign q[2] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40_combout ;

assign q[3] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53_combout ;

assign q[4] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66_combout ;

assign q[5] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79_combout ;

assign q[6] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92_combout ;

assign q[7] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105_combout ;

assign q[8] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118_combout ;

assign q[9] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131_combout ;

assign q[10] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144_combout ;

assign q[11] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157_combout ;

assign q[12] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170_combout ;

assign q[13] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183_combout ;

assign q[14] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196_combout ;

assign q[15] = \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209_combout ;

endmodule

module memory_LPM_RAM_DQ_1 (
	address_0,
	address_1,
	address_2,
	address_4,
	address_3,
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	data_0,
	we,
	data_1,
	data_2,
	data_3,
	data_4,
	data_5,
	data_6,
	data_7,
	data_8,
	data_9,
	data_10,
	data_11,
	data_12,
	data_13,
	data_14,
	data_15)/* synthesis synthesis_greybox=0 */;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_4;
input 	address_3;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
input 	data_0;
input 	we;
input 	data_1;
input 	data_2;
input 	data_3;
input 	data_4;
input 	data_5;
input 	data_6;
input 	data_7;
input 	data_8;
input 	data_9;
input 	data_10;
input 	data_11;
input 	data_12;
input 	data_13;
input 	data_14;
input 	data_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



memory_altram_1 sram(
	.address_0(address_0),
	.address_1(address_1),
	.address_2(address_2),
	.address_4(address_4),
	.address_3(address_3),
	.result_node_0(result_node_0),
	.result_node_1(result_node_1),
	.result_node_2(result_node_2),
	.result_node_3(result_node_3),
	.result_node_4(result_node_4),
	.result_node_5(result_node_5),
	.result_node_6(result_node_6),
	.result_node_7(result_node_7),
	.result_node_8(result_node_8),
	.result_node_9(result_node_9),
	.result_node_10(result_node_10),
	.result_node_11(result_node_11),
	.result_node_12(result_node_12),
	.result_node_13(result_node_13),
	.result_node_14(result_node_14),
	.result_node_15(result_node_15),
	.data_0(data_0),
	.we(we),
	.data_1(data_1),
	.data_2(data_2),
	.data_3(data_3),
	.data_4(data_4),
	.data_5(data_5),
	.data_6(data_6),
	.data_7(data_7),
	.data_8(data_8),
	.data_9(data_9),
	.data_10(data_10),
	.data_11(data_11),
	.data_12(data_12),
	.data_13(data_13),
	.data_14(data_14),
	.data_15(data_15));

endmodule

module memory_altram_1 (
	address_0,
	address_1,
	address_2,
	address_4,
	address_3,
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	data_0,
	we,
	data_1,
	data_2,
	data_3,
	data_4,
	data_5,
	data_6,
	data_7,
	data_8,
	data_9,
	data_10,
	data_11,
	data_12,
	data_13,
	data_14,
	data_15)/* synthesis synthesis_greybox=0 */;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_4;
input 	address_3;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
input 	data_0;
input 	we;
input 	data_1;
input 	data_2;
input 	data_3;
input 	data_4;
input 	data_5;
input 	data_6;
input 	data_7;
input 	data_8;
input 	data_9;
input 	data_10;
input 	data_11;
input 	data_12;
input 	data_13;
input 	data_14;
input 	data_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0_combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0_combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2_combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2_combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2_combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2_combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][0]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][1]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][2]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][3]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][4]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][5]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][6]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][7]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][8]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][9]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][10]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][11]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][12]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][13]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][14]~combout ;
wire \lpm_ram_dq_component|sram|latches[15][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[13][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[14][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[12][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[11][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[9][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[10][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[8][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[1][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[2][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[0][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[3][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[21][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[22][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[20][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[23][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[17][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[18][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[16][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[19][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[5][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[6][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[4][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[7][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[31][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[29][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[30][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[28][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[27][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[25][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[26][15]~combout ;
wire \lpm_ram_dq_component|sram|latches[24][15]~combout ;


memory_lpm_decode_1 decode(
	.address_0(address_0),
	.address_1(address_1),
	.address_2(address_2),
	.address_4(address_4),
	.address_3(address_3),
	.w_anode196w_2(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0_combout ),
	.w_anode287w_2(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0_combout ),
	.w_anode165w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2_combout ),
	.w_anode155w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2_combout ),
	.w_anode125w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2_combout ),
	.w_anode114w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2_combout ),
	.we(we),
	.w_anode135w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.w_anode43w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.w_anode16w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.w_anode226w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.w_anode205w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.w_anode317w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.w_anode185w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.w_anode165w_31(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.w_anode175w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.w_anode155w_31(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.w_anode145w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.w_anode125w_31(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.w_anode114w_31(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.w_anode33w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.w_anode53w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.w_anode256w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.w_anode266w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.w_anode246w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.w_anode276w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.w_anode216w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.w_anode236w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.w_anode73w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.w_anode83w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.w_anode63w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.w_anode93w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.w_anode367w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.w_anode347w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.w_anode357w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.w_anode337w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.w_anode327w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.w_anode307w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.w_anode296w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ));

memory_lpm_mux_1 mux(
	.address_0(address_0),
	.address_1(address_1),
	.address_2(address_2),
	.address_4(address_4),
	.address_3(address_3),
	.w_anode196w_2(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0_combout ),
	.w_anode287w_2(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0_combout ),
	.w_anode165w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2_combout ),
	.w_anode155w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2_combout ),
	.w_anode125w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2_combout ),
	.w_anode114w_3(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2_combout ),
	.result_node_0(result_node_0),
	.result_node_1(result_node_1),
	.result_node_2(result_node_2),
	.result_node_3(result_node_3),
	.result_node_4(result_node_4),
	.result_node_5(result_node_5),
	.result_node_6(result_node_6),
	.result_node_7(result_node_7),
	.result_node_8(result_node_8),
	.result_node_9(result_node_9),
	.result_node_10(result_node_10),
	.result_node_11(result_node_11),
	.result_node_12(result_node_12),
	.result_node_13(result_node_13),
	.result_node_14(result_node_14),
	.result_node_15(result_node_15),
	.latches_0_15(\lpm_ram_dq_component|sram|latches[15][0]~combout ),
	.latches_0_13(\lpm_ram_dq_component|sram|latches[13][0]~combout ),
	.latches_0_14(\lpm_ram_dq_component|sram|latches[14][0]~combout ),
	.latches_0_12(\lpm_ram_dq_component|sram|latches[12][0]~combout ),
	.latches_0_11(\lpm_ram_dq_component|sram|latches[11][0]~combout ),
	.latches_0_9(\lpm_ram_dq_component|sram|latches[9][0]~combout ),
	.latches_0_10(\lpm_ram_dq_component|sram|latches[10][0]~combout ),
	.latches_0_8(\lpm_ram_dq_component|sram|latches[8][0]~combout ),
	.latches_0_1(\lpm_ram_dq_component|sram|latches[1][0]~combout ),
	.latches_0_2(\lpm_ram_dq_component|sram|latches[2][0]~combout ),
	.latches_0_0(\lpm_ram_dq_component|sram|latches[0][0]~combout ),
	.latches_0_3(\lpm_ram_dq_component|sram|latches[3][0]~combout ),
	.latches_0_21(\lpm_ram_dq_component|sram|latches[21][0]~combout ),
	.latches_0_22(\lpm_ram_dq_component|sram|latches[22][0]~combout ),
	.latches_0_20(\lpm_ram_dq_component|sram|latches[20][0]~combout ),
	.latches_0_23(\lpm_ram_dq_component|sram|latches[23][0]~combout ),
	.latches_0_17(\lpm_ram_dq_component|sram|latches[17][0]~combout ),
	.latches_0_18(\lpm_ram_dq_component|sram|latches[18][0]~combout ),
	.latches_0_16(\lpm_ram_dq_component|sram|latches[16][0]~combout ),
	.latches_0_19(\lpm_ram_dq_component|sram|latches[19][0]~combout ),
	.latches_0_5(\lpm_ram_dq_component|sram|latches[5][0]~combout ),
	.latches_0_6(\lpm_ram_dq_component|sram|latches[6][0]~combout ),
	.latches_0_4(\lpm_ram_dq_component|sram|latches[4][0]~combout ),
	.latches_0_7(\lpm_ram_dq_component|sram|latches[7][0]~combout ),
	.latches_0_31(\lpm_ram_dq_component|sram|latches[31][0]~combout ),
	.latches_0_29(\lpm_ram_dq_component|sram|latches[29][0]~combout ),
	.latches_0_30(\lpm_ram_dq_component|sram|latches[30][0]~combout ),
	.latches_0_28(\lpm_ram_dq_component|sram|latches[28][0]~combout ),
	.latches_0_27(\lpm_ram_dq_component|sram|latches[27][0]~combout ),
	.latches_0_25(\lpm_ram_dq_component|sram|latches[25][0]~combout ),
	.latches_0_26(\lpm_ram_dq_component|sram|latches[26][0]~combout ),
	.latches_0_24(\lpm_ram_dq_component|sram|latches[24][0]~combout ),
	.latches_1_15(\lpm_ram_dq_component|sram|latches[15][1]~combout ),
	.latches_1_13(\lpm_ram_dq_component|sram|latches[13][1]~combout ),
	.latches_1_14(\lpm_ram_dq_component|sram|latches[14][1]~combout ),
	.latches_1_12(\lpm_ram_dq_component|sram|latches[12][1]~combout ),
	.latches_1_11(\lpm_ram_dq_component|sram|latches[11][1]~combout ),
	.latches_1_9(\lpm_ram_dq_component|sram|latches[9][1]~combout ),
	.latches_1_10(\lpm_ram_dq_component|sram|latches[10][1]~combout ),
	.latches_1_8(\lpm_ram_dq_component|sram|latches[8][1]~combout ),
	.latches_1_1(\lpm_ram_dq_component|sram|latches[1][1]~combout ),
	.latches_1_2(\lpm_ram_dq_component|sram|latches[2][1]~combout ),
	.latches_1_0(\lpm_ram_dq_component|sram|latches[0][1]~combout ),
	.latches_1_3(\lpm_ram_dq_component|sram|latches[3][1]~combout ),
	.latches_1_21(\lpm_ram_dq_component|sram|latches[21][1]~combout ),
	.latches_1_22(\lpm_ram_dq_component|sram|latches[22][1]~combout ),
	.latches_1_20(\lpm_ram_dq_component|sram|latches[20][1]~combout ),
	.latches_1_23(\lpm_ram_dq_component|sram|latches[23][1]~combout ),
	.latches_1_17(\lpm_ram_dq_component|sram|latches[17][1]~combout ),
	.latches_1_18(\lpm_ram_dq_component|sram|latches[18][1]~combout ),
	.latches_1_16(\lpm_ram_dq_component|sram|latches[16][1]~combout ),
	.latches_1_19(\lpm_ram_dq_component|sram|latches[19][1]~combout ),
	.latches_1_5(\lpm_ram_dq_component|sram|latches[5][1]~combout ),
	.latches_1_6(\lpm_ram_dq_component|sram|latches[6][1]~combout ),
	.latches_1_4(\lpm_ram_dq_component|sram|latches[4][1]~combout ),
	.latches_1_7(\lpm_ram_dq_component|sram|latches[7][1]~combout ),
	.latches_1_31(\lpm_ram_dq_component|sram|latches[31][1]~combout ),
	.latches_1_29(\lpm_ram_dq_component|sram|latches[29][1]~combout ),
	.latches_1_30(\lpm_ram_dq_component|sram|latches[30][1]~combout ),
	.latches_1_28(\lpm_ram_dq_component|sram|latches[28][1]~combout ),
	.latches_1_27(\lpm_ram_dq_component|sram|latches[27][1]~combout ),
	.latches_1_25(\lpm_ram_dq_component|sram|latches[25][1]~combout ),
	.latches_1_26(\lpm_ram_dq_component|sram|latches[26][1]~combout ),
	.latches_1_24(\lpm_ram_dq_component|sram|latches[24][1]~combout ),
	.latches_2_15(\lpm_ram_dq_component|sram|latches[15][2]~combout ),
	.latches_2_13(\lpm_ram_dq_component|sram|latches[13][2]~combout ),
	.latches_2_14(\lpm_ram_dq_component|sram|latches[14][2]~combout ),
	.latches_2_12(\lpm_ram_dq_component|sram|latches[12][2]~combout ),
	.latches_2_11(\lpm_ram_dq_component|sram|latches[11][2]~combout ),
	.latches_2_9(\lpm_ram_dq_component|sram|latches[9][2]~combout ),
	.latches_2_10(\lpm_ram_dq_component|sram|latches[10][2]~combout ),
	.latches_2_8(\lpm_ram_dq_component|sram|latches[8][2]~combout ),
	.latches_2_1(\lpm_ram_dq_component|sram|latches[1][2]~combout ),
	.latches_2_2(\lpm_ram_dq_component|sram|latches[2][2]~combout ),
	.latches_2_0(\lpm_ram_dq_component|sram|latches[0][2]~combout ),
	.latches_2_3(\lpm_ram_dq_component|sram|latches[3][2]~combout ),
	.latches_2_21(\lpm_ram_dq_component|sram|latches[21][2]~combout ),
	.latches_2_22(\lpm_ram_dq_component|sram|latches[22][2]~combout ),
	.latches_2_20(\lpm_ram_dq_component|sram|latches[20][2]~combout ),
	.latches_2_23(\lpm_ram_dq_component|sram|latches[23][2]~combout ),
	.latches_2_17(\lpm_ram_dq_component|sram|latches[17][2]~combout ),
	.latches_2_18(\lpm_ram_dq_component|sram|latches[18][2]~combout ),
	.latches_2_16(\lpm_ram_dq_component|sram|latches[16][2]~combout ),
	.latches_2_19(\lpm_ram_dq_component|sram|latches[19][2]~combout ),
	.latches_2_5(\lpm_ram_dq_component|sram|latches[5][2]~combout ),
	.latches_2_6(\lpm_ram_dq_component|sram|latches[6][2]~combout ),
	.latches_2_4(\lpm_ram_dq_component|sram|latches[4][2]~combout ),
	.latches_2_7(\lpm_ram_dq_component|sram|latches[7][2]~combout ),
	.latches_2_31(\lpm_ram_dq_component|sram|latches[31][2]~combout ),
	.latches_2_29(\lpm_ram_dq_component|sram|latches[29][2]~combout ),
	.latches_2_30(\lpm_ram_dq_component|sram|latches[30][2]~combout ),
	.latches_2_28(\lpm_ram_dq_component|sram|latches[28][2]~combout ),
	.latches_2_27(\lpm_ram_dq_component|sram|latches[27][2]~combout ),
	.latches_2_25(\lpm_ram_dq_component|sram|latches[25][2]~combout ),
	.latches_2_26(\lpm_ram_dq_component|sram|latches[26][2]~combout ),
	.latches_2_24(\lpm_ram_dq_component|sram|latches[24][2]~combout ),
	.latches_3_15(\lpm_ram_dq_component|sram|latches[15][3]~combout ),
	.latches_3_13(\lpm_ram_dq_component|sram|latches[13][3]~combout ),
	.latches_3_14(\lpm_ram_dq_component|sram|latches[14][3]~combout ),
	.latches_3_12(\lpm_ram_dq_component|sram|latches[12][3]~combout ),
	.latches_3_11(\lpm_ram_dq_component|sram|latches[11][3]~combout ),
	.latches_3_9(\lpm_ram_dq_component|sram|latches[9][3]~combout ),
	.latches_3_10(\lpm_ram_dq_component|sram|latches[10][3]~combout ),
	.latches_3_8(\lpm_ram_dq_component|sram|latches[8][3]~combout ),
	.latches_3_1(\lpm_ram_dq_component|sram|latches[1][3]~combout ),
	.latches_3_2(\lpm_ram_dq_component|sram|latches[2][3]~combout ),
	.latches_3_0(\lpm_ram_dq_component|sram|latches[0][3]~combout ),
	.latches_3_3(\lpm_ram_dq_component|sram|latches[3][3]~combout ),
	.latches_3_21(\lpm_ram_dq_component|sram|latches[21][3]~combout ),
	.latches_3_22(\lpm_ram_dq_component|sram|latches[22][3]~combout ),
	.latches_3_20(\lpm_ram_dq_component|sram|latches[20][3]~combout ),
	.latches_3_23(\lpm_ram_dq_component|sram|latches[23][3]~combout ),
	.latches_3_17(\lpm_ram_dq_component|sram|latches[17][3]~combout ),
	.latches_3_18(\lpm_ram_dq_component|sram|latches[18][3]~combout ),
	.latches_3_16(\lpm_ram_dq_component|sram|latches[16][3]~combout ),
	.latches_3_19(\lpm_ram_dq_component|sram|latches[19][3]~combout ),
	.latches_3_5(\lpm_ram_dq_component|sram|latches[5][3]~combout ),
	.latches_3_6(\lpm_ram_dq_component|sram|latches[6][3]~combout ),
	.latches_3_4(\lpm_ram_dq_component|sram|latches[4][3]~combout ),
	.latches_3_7(\lpm_ram_dq_component|sram|latches[7][3]~combout ),
	.latches_3_31(\lpm_ram_dq_component|sram|latches[31][3]~combout ),
	.latches_3_29(\lpm_ram_dq_component|sram|latches[29][3]~combout ),
	.latches_3_30(\lpm_ram_dq_component|sram|latches[30][3]~combout ),
	.latches_3_28(\lpm_ram_dq_component|sram|latches[28][3]~combout ),
	.latches_3_27(\lpm_ram_dq_component|sram|latches[27][3]~combout ),
	.latches_3_25(\lpm_ram_dq_component|sram|latches[25][3]~combout ),
	.latches_3_26(\lpm_ram_dq_component|sram|latches[26][3]~combout ),
	.latches_3_24(\lpm_ram_dq_component|sram|latches[24][3]~combout ),
	.latches_4_15(\lpm_ram_dq_component|sram|latches[15][4]~combout ),
	.latches_4_13(\lpm_ram_dq_component|sram|latches[13][4]~combout ),
	.latches_4_14(\lpm_ram_dq_component|sram|latches[14][4]~combout ),
	.latches_4_12(\lpm_ram_dq_component|sram|latches[12][4]~combout ),
	.latches_4_11(\lpm_ram_dq_component|sram|latches[11][4]~combout ),
	.latches_4_9(\lpm_ram_dq_component|sram|latches[9][4]~combout ),
	.latches_4_10(\lpm_ram_dq_component|sram|latches[10][4]~combout ),
	.latches_4_8(\lpm_ram_dq_component|sram|latches[8][4]~combout ),
	.latches_4_1(\lpm_ram_dq_component|sram|latches[1][4]~combout ),
	.latches_4_2(\lpm_ram_dq_component|sram|latches[2][4]~combout ),
	.latches_4_0(\lpm_ram_dq_component|sram|latches[0][4]~combout ),
	.latches_4_3(\lpm_ram_dq_component|sram|latches[3][4]~combout ),
	.latches_4_21(\lpm_ram_dq_component|sram|latches[21][4]~combout ),
	.latches_4_22(\lpm_ram_dq_component|sram|latches[22][4]~combout ),
	.latches_4_20(\lpm_ram_dq_component|sram|latches[20][4]~combout ),
	.latches_4_23(\lpm_ram_dq_component|sram|latches[23][4]~combout ),
	.latches_4_17(\lpm_ram_dq_component|sram|latches[17][4]~combout ),
	.latches_4_18(\lpm_ram_dq_component|sram|latches[18][4]~combout ),
	.latches_4_16(\lpm_ram_dq_component|sram|latches[16][4]~combout ),
	.latches_4_19(\lpm_ram_dq_component|sram|latches[19][4]~combout ),
	.latches_4_5(\lpm_ram_dq_component|sram|latches[5][4]~combout ),
	.latches_4_6(\lpm_ram_dq_component|sram|latches[6][4]~combout ),
	.latches_4_4(\lpm_ram_dq_component|sram|latches[4][4]~combout ),
	.latches_4_7(\lpm_ram_dq_component|sram|latches[7][4]~combout ),
	.latches_4_31(\lpm_ram_dq_component|sram|latches[31][4]~combout ),
	.latches_4_29(\lpm_ram_dq_component|sram|latches[29][4]~combout ),
	.latches_4_30(\lpm_ram_dq_component|sram|latches[30][4]~combout ),
	.latches_4_28(\lpm_ram_dq_component|sram|latches[28][4]~combout ),
	.latches_4_27(\lpm_ram_dq_component|sram|latches[27][4]~combout ),
	.latches_4_25(\lpm_ram_dq_component|sram|latches[25][4]~combout ),
	.latches_4_26(\lpm_ram_dq_component|sram|latches[26][4]~combout ),
	.latches_4_24(\lpm_ram_dq_component|sram|latches[24][4]~combout ),
	.latches_5_15(\lpm_ram_dq_component|sram|latches[15][5]~combout ),
	.latches_5_13(\lpm_ram_dq_component|sram|latches[13][5]~combout ),
	.latches_5_14(\lpm_ram_dq_component|sram|latches[14][5]~combout ),
	.latches_5_12(\lpm_ram_dq_component|sram|latches[12][5]~combout ),
	.latches_5_11(\lpm_ram_dq_component|sram|latches[11][5]~combout ),
	.latches_5_9(\lpm_ram_dq_component|sram|latches[9][5]~combout ),
	.latches_5_10(\lpm_ram_dq_component|sram|latches[10][5]~combout ),
	.latches_5_8(\lpm_ram_dq_component|sram|latches[8][5]~combout ),
	.latches_5_1(\lpm_ram_dq_component|sram|latches[1][5]~combout ),
	.latches_5_2(\lpm_ram_dq_component|sram|latches[2][5]~combout ),
	.latches_5_0(\lpm_ram_dq_component|sram|latches[0][5]~combout ),
	.latches_5_3(\lpm_ram_dq_component|sram|latches[3][5]~combout ),
	.latches_5_21(\lpm_ram_dq_component|sram|latches[21][5]~combout ),
	.latches_5_22(\lpm_ram_dq_component|sram|latches[22][5]~combout ),
	.latches_5_20(\lpm_ram_dq_component|sram|latches[20][5]~combout ),
	.latches_5_23(\lpm_ram_dq_component|sram|latches[23][5]~combout ),
	.latches_5_17(\lpm_ram_dq_component|sram|latches[17][5]~combout ),
	.latches_5_18(\lpm_ram_dq_component|sram|latches[18][5]~combout ),
	.latches_5_16(\lpm_ram_dq_component|sram|latches[16][5]~combout ),
	.latches_5_19(\lpm_ram_dq_component|sram|latches[19][5]~combout ),
	.latches_5_5(\lpm_ram_dq_component|sram|latches[5][5]~combout ),
	.latches_5_6(\lpm_ram_dq_component|sram|latches[6][5]~combout ),
	.latches_5_4(\lpm_ram_dq_component|sram|latches[4][5]~combout ),
	.latches_5_7(\lpm_ram_dq_component|sram|latches[7][5]~combout ),
	.latches_5_31(\lpm_ram_dq_component|sram|latches[31][5]~combout ),
	.latches_5_29(\lpm_ram_dq_component|sram|latches[29][5]~combout ),
	.latches_5_30(\lpm_ram_dq_component|sram|latches[30][5]~combout ),
	.latches_5_28(\lpm_ram_dq_component|sram|latches[28][5]~combout ),
	.latches_5_27(\lpm_ram_dq_component|sram|latches[27][5]~combout ),
	.latches_5_25(\lpm_ram_dq_component|sram|latches[25][5]~combout ),
	.latches_5_26(\lpm_ram_dq_component|sram|latches[26][5]~combout ),
	.latches_5_24(\lpm_ram_dq_component|sram|latches[24][5]~combout ),
	.latches_6_15(\lpm_ram_dq_component|sram|latches[15][6]~combout ),
	.latches_6_13(\lpm_ram_dq_component|sram|latches[13][6]~combout ),
	.latches_6_14(\lpm_ram_dq_component|sram|latches[14][6]~combout ),
	.latches_6_12(\lpm_ram_dq_component|sram|latches[12][6]~combout ),
	.latches_6_11(\lpm_ram_dq_component|sram|latches[11][6]~combout ),
	.latches_6_9(\lpm_ram_dq_component|sram|latches[9][6]~combout ),
	.latches_6_10(\lpm_ram_dq_component|sram|latches[10][6]~combout ),
	.latches_6_8(\lpm_ram_dq_component|sram|latches[8][6]~combout ),
	.latches_6_1(\lpm_ram_dq_component|sram|latches[1][6]~combout ),
	.latches_6_2(\lpm_ram_dq_component|sram|latches[2][6]~combout ),
	.latches_6_0(\lpm_ram_dq_component|sram|latches[0][6]~combout ),
	.latches_6_3(\lpm_ram_dq_component|sram|latches[3][6]~combout ),
	.latches_6_21(\lpm_ram_dq_component|sram|latches[21][6]~combout ),
	.latches_6_22(\lpm_ram_dq_component|sram|latches[22][6]~combout ),
	.latches_6_20(\lpm_ram_dq_component|sram|latches[20][6]~combout ),
	.latches_6_23(\lpm_ram_dq_component|sram|latches[23][6]~combout ),
	.latches_6_17(\lpm_ram_dq_component|sram|latches[17][6]~combout ),
	.latches_6_18(\lpm_ram_dq_component|sram|latches[18][6]~combout ),
	.latches_6_16(\lpm_ram_dq_component|sram|latches[16][6]~combout ),
	.latches_6_19(\lpm_ram_dq_component|sram|latches[19][6]~combout ),
	.latches_6_5(\lpm_ram_dq_component|sram|latches[5][6]~combout ),
	.latches_6_6(\lpm_ram_dq_component|sram|latches[6][6]~combout ),
	.latches_6_4(\lpm_ram_dq_component|sram|latches[4][6]~combout ),
	.latches_6_7(\lpm_ram_dq_component|sram|latches[7][6]~combout ),
	.latches_6_31(\lpm_ram_dq_component|sram|latches[31][6]~combout ),
	.latches_6_29(\lpm_ram_dq_component|sram|latches[29][6]~combout ),
	.latches_6_30(\lpm_ram_dq_component|sram|latches[30][6]~combout ),
	.latches_6_28(\lpm_ram_dq_component|sram|latches[28][6]~combout ),
	.latches_6_27(\lpm_ram_dq_component|sram|latches[27][6]~combout ),
	.latches_6_25(\lpm_ram_dq_component|sram|latches[25][6]~combout ),
	.latches_6_26(\lpm_ram_dq_component|sram|latches[26][6]~combout ),
	.latches_6_24(\lpm_ram_dq_component|sram|latches[24][6]~combout ),
	.latches_7_15(\lpm_ram_dq_component|sram|latches[15][7]~combout ),
	.latches_7_13(\lpm_ram_dq_component|sram|latches[13][7]~combout ),
	.latches_7_14(\lpm_ram_dq_component|sram|latches[14][7]~combout ),
	.latches_7_12(\lpm_ram_dq_component|sram|latches[12][7]~combout ),
	.latches_7_11(\lpm_ram_dq_component|sram|latches[11][7]~combout ),
	.latches_7_9(\lpm_ram_dq_component|sram|latches[9][7]~combout ),
	.latches_7_10(\lpm_ram_dq_component|sram|latches[10][7]~combout ),
	.latches_7_8(\lpm_ram_dq_component|sram|latches[8][7]~combout ),
	.latches_7_1(\lpm_ram_dq_component|sram|latches[1][7]~combout ),
	.latches_7_2(\lpm_ram_dq_component|sram|latches[2][7]~combout ),
	.latches_7_0(\lpm_ram_dq_component|sram|latches[0][7]~combout ),
	.latches_7_3(\lpm_ram_dq_component|sram|latches[3][7]~combout ),
	.latches_7_21(\lpm_ram_dq_component|sram|latches[21][7]~combout ),
	.latches_7_22(\lpm_ram_dq_component|sram|latches[22][7]~combout ),
	.latches_7_20(\lpm_ram_dq_component|sram|latches[20][7]~combout ),
	.latches_7_23(\lpm_ram_dq_component|sram|latches[23][7]~combout ),
	.latches_7_17(\lpm_ram_dq_component|sram|latches[17][7]~combout ),
	.latches_7_18(\lpm_ram_dq_component|sram|latches[18][7]~combout ),
	.latches_7_16(\lpm_ram_dq_component|sram|latches[16][7]~combout ),
	.latches_7_19(\lpm_ram_dq_component|sram|latches[19][7]~combout ),
	.latches_7_5(\lpm_ram_dq_component|sram|latches[5][7]~combout ),
	.latches_7_6(\lpm_ram_dq_component|sram|latches[6][7]~combout ),
	.latches_7_4(\lpm_ram_dq_component|sram|latches[4][7]~combout ),
	.latches_7_7(\lpm_ram_dq_component|sram|latches[7][7]~combout ),
	.latches_7_31(\lpm_ram_dq_component|sram|latches[31][7]~combout ),
	.latches_7_29(\lpm_ram_dq_component|sram|latches[29][7]~combout ),
	.latches_7_30(\lpm_ram_dq_component|sram|latches[30][7]~combout ),
	.latches_7_28(\lpm_ram_dq_component|sram|latches[28][7]~combout ),
	.latches_7_27(\lpm_ram_dq_component|sram|latches[27][7]~combout ),
	.latches_7_25(\lpm_ram_dq_component|sram|latches[25][7]~combout ),
	.latches_7_26(\lpm_ram_dq_component|sram|latches[26][7]~combout ),
	.latches_7_24(\lpm_ram_dq_component|sram|latches[24][7]~combout ),
	.latches_8_15(\lpm_ram_dq_component|sram|latches[15][8]~combout ),
	.latches_8_13(\lpm_ram_dq_component|sram|latches[13][8]~combout ),
	.latches_8_14(\lpm_ram_dq_component|sram|latches[14][8]~combout ),
	.latches_8_12(\lpm_ram_dq_component|sram|latches[12][8]~combout ),
	.latches_8_11(\lpm_ram_dq_component|sram|latches[11][8]~combout ),
	.latches_8_9(\lpm_ram_dq_component|sram|latches[9][8]~combout ),
	.latches_8_10(\lpm_ram_dq_component|sram|latches[10][8]~combout ),
	.latches_8_8(\lpm_ram_dq_component|sram|latches[8][8]~combout ),
	.latches_8_1(\lpm_ram_dq_component|sram|latches[1][8]~combout ),
	.latches_8_2(\lpm_ram_dq_component|sram|latches[2][8]~combout ),
	.latches_8_0(\lpm_ram_dq_component|sram|latches[0][8]~combout ),
	.latches_8_3(\lpm_ram_dq_component|sram|latches[3][8]~combout ),
	.latches_8_21(\lpm_ram_dq_component|sram|latches[21][8]~combout ),
	.latches_8_22(\lpm_ram_dq_component|sram|latches[22][8]~combout ),
	.latches_8_20(\lpm_ram_dq_component|sram|latches[20][8]~combout ),
	.latches_8_23(\lpm_ram_dq_component|sram|latches[23][8]~combout ),
	.latches_8_17(\lpm_ram_dq_component|sram|latches[17][8]~combout ),
	.latches_8_18(\lpm_ram_dq_component|sram|latches[18][8]~combout ),
	.latches_8_16(\lpm_ram_dq_component|sram|latches[16][8]~combout ),
	.latches_8_19(\lpm_ram_dq_component|sram|latches[19][8]~combout ),
	.latches_8_5(\lpm_ram_dq_component|sram|latches[5][8]~combout ),
	.latches_8_6(\lpm_ram_dq_component|sram|latches[6][8]~combout ),
	.latches_8_4(\lpm_ram_dq_component|sram|latches[4][8]~combout ),
	.latches_8_7(\lpm_ram_dq_component|sram|latches[7][8]~combout ),
	.latches_8_31(\lpm_ram_dq_component|sram|latches[31][8]~combout ),
	.latches_8_29(\lpm_ram_dq_component|sram|latches[29][8]~combout ),
	.latches_8_30(\lpm_ram_dq_component|sram|latches[30][8]~combout ),
	.latches_8_28(\lpm_ram_dq_component|sram|latches[28][8]~combout ),
	.latches_8_27(\lpm_ram_dq_component|sram|latches[27][8]~combout ),
	.latches_8_25(\lpm_ram_dq_component|sram|latches[25][8]~combout ),
	.latches_8_26(\lpm_ram_dq_component|sram|latches[26][8]~combout ),
	.latches_8_24(\lpm_ram_dq_component|sram|latches[24][8]~combout ),
	.latches_9_15(\lpm_ram_dq_component|sram|latches[15][9]~combout ),
	.latches_9_13(\lpm_ram_dq_component|sram|latches[13][9]~combout ),
	.latches_9_14(\lpm_ram_dq_component|sram|latches[14][9]~combout ),
	.latches_9_12(\lpm_ram_dq_component|sram|latches[12][9]~combout ),
	.latches_9_11(\lpm_ram_dq_component|sram|latches[11][9]~combout ),
	.latches_9_9(\lpm_ram_dq_component|sram|latches[9][9]~combout ),
	.latches_9_10(\lpm_ram_dq_component|sram|latches[10][9]~combout ),
	.latches_9_8(\lpm_ram_dq_component|sram|latches[8][9]~combout ),
	.latches_9_1(\lpm_ram_dq_component|sram|latches[1][9]~combout ),
	.latches_9_2(\lpm_ram_dq_component|sram|latches[2][9]~combout ),
	.latches_9_0(\lpm_ram_dq_component|sram|latches[0][9]~combout ),
	.latches_9_3(\lpm_ram_dq_component|sram|latches[3][9]~combout ),
	.latches_9_21(\lpm_ram_dq_component|sram|latches[21][9]~combout ),
	.latches_9_22(\lpm_ram_dq_component|sram|latches[22][9]~combout ),
	.latches_9_20(\lpm_ram_dq_component|sram|latches[20][9]~combout ),
	.latches_9_23(\lpm_ram_dq_component|sram|latches[23][9]~combout ),
	.latches_9_17(\lpm_ram_dq_component|sram|latches[17][9]~combout ),
	.latches_9_18(\lpm_ram_dq_component|sram|latches[18][9]~combout ),
	.latches_9_16(\lpm_ram_dq_component|sram|latches[16][9]~combout ),
	.latches_9_19(\lpm_ram_dq_component|sram|latches[19][9]~combout ),
	.latches_9_5(\lpm_ram_dq_component|sram|latches[5][9]~combout ),
	.latches_9_6(\lpm_ram_dq_component|sram|latches[6][9]~combout ),
	.latches_9_4(\lpm_ram_dq_component|sram|latches[4][9]~combout ),
	.latches_9_7(\lpm_ram_dq_component|sram|latches[7][9]~combout ),
	.latches_9_31(\lpm_ram_dq_component|sram|latches[31][9]~combout ),
	.latches_9_29(\lpm_ram_dq_component|sram|latches[29][9]~combout ),
	.latches_9_30(\lpm_ram_dq_component|sram|latches[30][9]~combout ),
	.latches_9_28(\lpm_ram_dq_component|sram|latches[28][9]~combout ),
	.latches_9_27(\lpm_ram_dq_component|sram|latches[27][9]~combout ),
	.latches_9_25(\lpm_ram_dq_component|sram|latches[25][9]~combout ),
	.latches_9_26(\lpm_ram_dq_component|sram|latches[26][9]~combout ),
	.latches_9_24(\lpm_ram_dq_component|sram|latches[24][9]~combout ),
	.latches_10_15(\lpm_ram_dq_component|sram|latches[15][10]~combout ),
	.latches_10_13(\lpm_ram_dq_component|sram|latches[13][10]~combout ),
	.latches_10_14(\lpm_ram_dq_component|sram|latches[14][10]~combout ),
	.latches_10_12(\lpm_ram_dq_component|sram|latches[12][10]~combout ),
	.latches_10_11(\lpm_ram_dq_component|sram|latches[11][10]~combout ),
	.latches_10_9(\lpm_ram_dq_component|sram|latches[9][10]~combout ),
	.latches_10_10(\lpm_ram_dq_component|sram|latches[10][10]~combout ),
	.latches_10_8(\lpm_ram_dq_component|sram|latches[8][10]~combout ),
	.latches_10_1(\lpm_ram_dq_component|sram|latches[1][10]~combout ),
	.latches_10_2(\lpm_ram_dq_component|sram|latches[2][10]~combout ),
	.latches_10_0(\lpm_ram_dq_component|sram|latches[0][10]~combout ),
	.latches_10_3(\lpm_ram_dq_component|sram|latches[3][10]~combout ),
	.latches_10_21(\lpm_ram_dq_component|sram|latches[21][10]~combout ),
	.latches_10_22(\lpm_ram_dq_component|sram|latches[22][10]~combout ),
	.latches_10_20(\lpm_ram_dq_component|sram|latches[20][10]~combout ),
	.latches_10_23(\lpm_ram_dq_component|sram|latches[23][10]~combout ),
	.latches_10_17(\lpm_ram_dq_component|sram|latches[17][10]~combout ),
	.latches_10_18(\lpm_ram_dq_component|sram|latches[18][10]~combout ),
	.latches_10_16(\lpm_ram_dq_component|sram|latches[16][10]~combout ),
	.latches_10_19(\lpm_ram_dq_component|sram|latches[19][10]~combout ),
	.latches_10_5(\lpm_ram_dq_component|sram|latches[5][10]~combout ),
	.latches_10_6(\lpm_ram_dq_component|sram|latches[6][10]~combout ),
	.latches_10_4(\lpm_ram_dq_component|sram|latches[4][10]~combout ),
	.latches_10_7(\lpm_ram_dq_component|sram|latches[7][10]~combout ),
	.latches_10_31(\lpm_ram_dq_component|sram|latches[31][10]~combout ),
	.latches_10_29(\lpm_ram_dq_component|sram|latches[29][10]~combout ),
	.latches_10_30(\lpm_ram_dq_component|sram|latches[30][10]~combout ),
	.latches_10_28(\lpm_ram_dq_component|sram|latches[28][10]~combout ),
	.latches_10_27(\lpm_ram_dq_component|sram|latches[27][10]~combout ),
	.latches_10_25(\lpm_ram_dq_component|sram|latches[25][10]~combout ),
	.latches_10_26(\lpm_ram_dq_component|sram|latches[26][10]~combout ),
	.latches_10_24(\lpm_ram_dq_component|sram|latches[24][10]~combout ),
	.latches_11_15(\lpm_ram_dq_component|sram|latches[15][11]~combout ),
	.latches_11_13(\lpm_ram_dq_component|sram|latches[13][11]~combout ),
	.latches_11_14(\lpm_ram_dq_component|sram|latches[14][11]~combout ),
	.latches_11_12(\lpm_ram_dq_component|sram|latches[12][11]~combout ),
	.latches_11_11(\lpm_ram_dq_component|sram|latches[11][11]~combout ),
	.latches_11_9(\lpm_ram_dq_component|sram|latches[9][11]~combout ),
	.latches_11_10(\lpm_ram_dq_component|sram|latches[10][11]~combout ),
	.latches_11_8(\lpm_ram_dq_component|sram|latches[8][11]~combout ),
	.latches_11_1(\lpm_ram_dq_component|sram|latches[1][11]~combout ),
	.latches_11_2(\lpm_ram_dq_component|sram|latches[2][11]~combout ),
	.latches_11_0(\lpm_ram_dq_component|sram|latches[0][11]~combout ),
	.latches_11_3(\lpm_ram_dq_component|sram|latches[3][11]~combout ),
	.latches_11_21(\lpm_ram_dq_component|sram|latches[21][11]~combout ),
	.latches_11_22(\lpm_ram_dq_component|sram|latches[22][11]~combout ),
	.latches_11_20(\lpm_ram_dq_component|sram|latches[20][11]~combout ),
	.latches_11_23(\lpm_ram_dq_component|sram|latches[23][11]~combout ),
	.latches_11_17(\lpm_ram_dq_component|sram|latches[17][11]~combout ),
	.latches_11_18(\lpm_ram_dq_component|sram|latches[18][11]~combout ),
	.latches_11_16(\lpm_ram_dq_component|sram|latches[16][11]~combout ),
	.latches_11_19(\lpm_ram_dq_component|sram|latches[19][11]~combout ),
	.latches_11_5(\lpm_ram_dq_component|sram|latches[5][11]~combout ),
	.latches_11_6(\lpm_ram_dq_component|sram|latches[6][11]~combout ),
	.latches_11_4(\lpm_ram_dq_component|sram|latches[4][11]~combout ),
	.latches_11_7(\lpm_ram_dq_component|sram|latches[7][11]~combout ),
	.latches_11_31(\lpm_ram_dq_component|sram|latches[31][11]~combout ),
	.latches_11_29(\lpm_ram_dq_component|sram|latches[29][11]~combout ),
	.latches_11_30(\lpm_ram_dq_component|sram|latches[30][11]~combout ),
	.latches_11_28(\lpm_ram_dq_component|sram|latches[28][11]~combout ),
	.latches_11_27(\lpm_ram_dq_component|sram|latches[27][11]~combout ),
	.latches_11_25(\lpm_ram_dq_component|sram|latches[25][11]~combout ),
	.latches_11_26(\lpm_ram_dq_component|sram|latches[26][11]~combout ),
	.latches_11_24(\lpm_ram_dq_component|sram|latches[24][11]~combout ),
	.latches_12_15(\lpm_ram_dq_component|sram|latches[15][12]~combout ),
	.latches_12_13(\lpm_ram_dq_component|sram|latches[13][12]~combout ),
	.latches_12_14(\lpm_ram_dq_component|sram|latches[14][12]~combout ),
	.latches_12_12(\lpm_ram_dq_component|sram|latches[12][12]~combout ),
	.latches_12_11(\lpm_ram_dq_component|sram|latches[11][12]~combout ),
	.latches_12_9(\lpm_ram_dq_component|sram|latches[9][12]~combout ),
	.latches_12_10(\lpm_ram_dq_component|sram|latches[10][12]~combout ),
	.latches_12_8(\lpm_ram_dq_component|sram|latches[8][12]~combout ),
	.latches_12_1(\lpm_ram_dq_component|sram|latches[1][12]~combout ),
	.latches_12_2(\lpm_ram_dq_component|sram|latches[2][12]~combout ),
	.latches_12_0(\lpm_ram_dq_component|sram|latches[0][12]~combout ),
	.latches_12_3(\lpm_ram_dq_component|sram|latches[3][12]~combout ),
	.latches_12_21(\lpm_ram_dq_component|sram|latches[21][12]~combout ),
	.latches_12_22(\lpm_ram_dq_component|sram|latches[22][12]~combout ),
	.latches_12_20(\lpm_ram_dq_component|sram|latches[20][12]~combout ),
	.latches_12_23(\lpm_ram_dq_component|sram|latches[23][12]~combout ),
	.latches_12_17(\lpm_ram_dq_component|sram|latches[17][12]~combout ),
	.latches_12_18(\lpm_ram_dq_component|sram|latches[18][12]~combout ),
	.latches_12_16(\lpm_ram_dq_component|sram|latches[16][12]~combout ),
	.latches_12_19(\lpm_ram_dq_component|sram|latches[19][12]~combout ),
	.latches_12_5(\lpm_ram_dq_component|sram|latches[5][12]~combout ),
	.latches_12_6(\lpm_ram_dq_component|sram|latches[6][12]~combout ),
	.latches_12_4(\lpm_ram_dq_component|sram|latches[4][12]~combout ),
	.latches_12_7(\lpm_ram_dq_component|sram|latches[7][12]~combout ),
	.latches_12_31(\lpm_ram_dq_component|sram|latches[31][12]~combout ),
	.latches_12_29(\lpm_ram_dq_component|sram|latches[29][12]~combout ),
	.latches_12_30(\lpm_ram_dq_component|sram|latches[30][12]~combout ),
	.latches_12_28(\lpm_ram_dq_component|sram|latches[28][12]~combout ),
	.latches_12_27(\lpm_ram_dq_component|sram|latches[27][12]~combout ),
	.latches_12_25(\lpm_ram_dq_component|sram|latches[25][12]~combout ),
	.latches_12_26(\lpm_ram_dq_component|sram|latches[26][12]~combout ),
	.latches_12_24(\lpm_ram_dq_component|sram|latches[24][12]~combout ),
	.latches_13_15(\lpm_ram_dq_component|sram|latches[15][13]~combout ),
	.latches_13_13(\lpm_ram_dq_component|sram|latches[13][13]~combout ),
	.latches_13_14(\lpm_ram_dq_component|sram|latches[14][13]~combout ),
	.latches_13_12(\lpm_ram_dq_component|sram|latches[12][13]~combout ),
	.latches_13_11(\lpm_ram_dq_component|sram|latches[11][13]~combout ),
	.latches_13_9(\lpm_ram_dq_component|sram|latches[9][13]~combout ),
	.latches_13_10(\lpm_ram_dq_component|sram|latches[10][13]~combout ),
	.latches_13_8(\lpm_ram_dq_component|sram|latches[8][13]~combout ),
	.latches_13_1(\lpm_ram_dq_component|sram|latches[1][13]~combout ),
	.latches_13_2(\lpm_ram_dq_component|sram|latches[2][13]~combout ),
	.latches_13_0(\lpm_ram_dq_component|sram|latches[0][13]~combout ),
	.latches_13_3(\lpm_ram_dq_component|sram|latches[3][13]~combout ),
	.latches_13_21(\lpm_ram_dq_component|sram|latches[21][13]~combout ),
	.latches_13_22(\lpm_ram_dq_component|sram|latches[22][13]~combout ),
	.latches_13_20(\lpm_ram_dq_component|sram|latches[20][13]~combout ),
	.latches_13_23(\lpm_ram_dq_component|sram|latches[23][13]~combout ),
	.latches_13_17(\lpm_ram_dq_component|sram|latches[17][13]~combout ),
	.latches_13_18(\lpm_ram_dq_component|sram|latches[18][13]~combout ),
	.latches_13_16(\lpm_ram_dq_component|sram|latches[16][13]~combout ),
	.latches_13_19(\lpm_ram_dq_component|sram|latches[19][13]~combout ),
	.latches_13_5(\lpm_ram_dq_component|sram|latches[5][13]~combout ),
	.latches_13_6(\lpm_ram_dq_component|sram|latches[6][13]~combout ),
	.latches_13_4(\lpm_ram_dq_component|sram|latches[4][13]~combout ),
	.latches_13_7(\lpm_ram_dq_component|sram|latches[7][13]~combout ),
	.latches_13_31(\lpm_ram_dq_component|sram|latches[31][13]~combout ),
	.latches_13_29(\lpm_ram_dq_component|sram|latches[29][13]~combout ),
	.latches_13_30(\lpm_ram_dq_component|sram|latches[30][13]~combout ),
	.latches_13_28(\lpm_ram_dq_component|sram|latches[28][13]~combout ),
	.latches_13_27(\lpm_ram_dq_component|sram|latches[27][13]~combout ),
	.latches_13_25(\lpm_ram_dq_component|sram|latches[25][13]~combout ),
	.latches_13_26(\lpm_ram_dq_component|sram|latches[26][13]~combout ),
	.latches_13_24(\lpm_ram_dq_component|sram|latches[24][13]~combout ),
	.latches_14_15(\lpm_ram_dq_component|sram|latches[15][14]~combout ),
	.latches_14_13(\lpm_ram_dq_component|sram|latches[13][14]~combout ),
	.latches_14_14(\lpm_ram_dq_component|sram|latches[14][14]~combout ),
	.latches_14_12(\lpm_ram_dq_component|sram|latches[12][14]~combout ),
	.latches_14_11(\lpm_ram_dq_component|sram|latches[11][14]~combout ),
	.latches_14_9(\lpm_ram_dq_component|sram|latches[9][14]~combout ),
	.latches_14_10(\lpm_ram_dq_component|sram|latches[10][14]~combout ),
	.latches_14_8(\lpm_ram_dq_component|sram|latches[8][14]~combout ),
	.latches_14_1(\lpm_ram_dq_component|sram|latches[1][14]~combout ),
	.latches_14_2(\lpm_ram_dq_component|sram|latches[2][14]~combout ),
	.latches_14_0(\lpm_ram_dq_component|sram|latches[0][14]~combout ),
	.latches_14_3(\lpm_ram_dq_component|sram|latches[3][14]~combout ),
	.latches_14_21(\lpm_ram_dq_component|sram|latches[21][14]~combout ),
	.latches_14_22(\lpm_ram_dq_component|sram|latches[22][14]~combout ),
	.latches_14_20(\lpm_ram_dq_component|sram|latches[20][14]~combout ),
	.latches_14_23(\lpm_ram_dq_component|sram|latches[23][14]~combout ),
	.latches_14_17(\lpm_ram_dq_component|sram|latches[17][14]~combout ),
	.latches_14_18(\lpm_ram_dq_component|sram|latches[18][14]~combout ),
	.latches_14_16(\lpm_ram_dq_component|sram|latches[16][14]~combout ),
	.latches_14_19(\lpm_ram_dq_component|sram|latches[19][14]~combout ),
	.latches_14_5(\lpm_ram_dq_component|sram|latches[5][14]~combout ),
	.latches_14_6(\lpm_ram_dq_component|sram|latches[6][14]~combout ),
	.latches_14_4(\lpm_ram_dq_component|sram|latches[4][14]~combout ),
	.latches_14_7(\lpm_ram_dq_component|sram|latches[7][14]~combout ),
	.latches_14_31(\lpm_ram_dq_component|sram|latches[31][14]~combout ),
	.latches_14_29(\lpm_ram_dq_component|sram|latches[29][14]~combout ),
	.latches_14_30(\lpm_ram_dq_component|sram|latches[30][14]~combout ),
	.latches_14_28(\lpm_ram_dq_component|sram|latches[28][14]~combout ),
	.latches_14_27(\lpm_ram_dq_component|sram|latches[27][14]~combout ),
	.latches_14_25(\lpm_ram_dq_component|sram|latches[25][14]~combout ),
	.latches_14_26(\lpm_ram_dq_component|sram|latches[26][14]~combout ),
	.latches_14_24(\lpm_ram_dq_component|sram|latches[24][14]~combout ),
	.latches_15_15(\lpm_ram_dq_component|sram|latches[15][15]~combout ),
	.latches_15_13(\lpm_ram_dq_component|sram|latches[13][15]~combout ),
	.latches_15_14(\lpm_ram_dq_component|sram|latches[14][15]~combout ),
	.latches_15_12(\lpm_ram_dq_component|sram|latches[12][15]~combout ),
	.latches_15_11(\lpm_ram_dq_component|sram|latches[11][15]~combout ),
	.latches_15_9(\lpm_ram_dq_component|sram|latches[9][15]~combout ),
	.latches_15_10(\lpm_ram_dq_component|sram|latches[10][15]~combout ),
	.latches_15_8(\lpm_ram_dq_component|sram|latches[8][15]~combout ),
	.latches_15_1(\lpm_ram_dq_component|sram|latches[1][15]~combout ),
	.latches_15_2(\lpm_ram_dq_component|sram|latches[2][15]~combout ),
	.latches_15_0(\lpm_ram_dq_component|sram|latches[0][15]~combout ),
	.latches_15_3(\lpm_ram_dq_component|sram|latches[3][15]~combout ),
	.latches_15_21(\lpm_ram_dq_component|sram|latches[21][15]~combout ),
	.latches_15_22(\lpm_ram_dq_component|sram|latches[22][15]~combout ),
	.latches_15_20(\lpm_ram_dq_component|sram|latches[20][15]~combout ),
	.latches_15_23(\lpm_ram_dq_component|sram|latches[23][15]~combout ),
	.latches_15_17(\lpm_ram_dq_component|sram|latches[17][15]~combout ),
	.latches_15_18(\lpm_ram_dq_component|sram|latches[18][15]~combout ),
	.latches_15_16(\lpm_ram_dq_component|sram|latches[16][15]~combout ),
	.latches_15_19(\lpm_ram_dq_component|sram|latches[19][15]~combout ),
	.latches_15_5(\lpm_ram_dq_component|sram|latches[5][15]~combout ),
	.latches_15_6(\lpm_ram_dq_component|sram|latches[6][15]~combout ),
	.latches_15_4(\lpm_ram_dq_component|sram|latches[4][15]~combout ),
	.latches_15_7(\lpm_ram_dq_component|sram|latches[7][15]~combout ),
	.latches_15_31(\lpm_ram_dq_component|sram|latches[31][15]~combout ),
	.latches_15_29(\lpm_ram_dq_component|sram|latches[29][15]~combout ),
	.latches_15_30(\lpm_ram_dq_component|sram|latches[30][15]~combout ),
	.latches_15_28(\lpm_ram_dq_component|sram|latches[28][15]~combout ),
	.latches_15_27(\lpm_ram_dq_component|sram|latches[27][15]~combout ),
	.latches_15_25(\lpm_ram_dq_component|sram|latches[25][15]~combout ),
	.latches_15_26(\lpm_ram_dq_component|sram|latches[26][15]~combout ),
	.latches_15_24(\lpm_ram_dq_component|sram|latches[24][15]~combout ));

maxv_lcell \lpm_ram_dq_component|sram|latches[15][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[15][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[13][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[14][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[12][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[11][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[9][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[10][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[8][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[1][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[2][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[0][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[3][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[21][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[22][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[20][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[23][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[17][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[18][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[16][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[19][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[5][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[6][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[4][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[7][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[31][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[29][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[30][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[28][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[27][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[25][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[26][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][0] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_0),
	.datac(\lpm_ram_dq_component|sram|latches[24][0]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][0]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][0] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][0] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][0] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][0] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][0] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][0] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[15][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[13][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[14][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[12][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[11][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[9][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[10][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[8][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[1][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[2][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[0][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[3][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[21][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[22][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[20][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[23][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[17][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[18][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[16][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[19][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[5][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[6][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[4][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[7][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[31][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[29][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[30][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[28][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[27][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[25][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[26][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][1] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_1),
	.datac(\lpm_ram_dq_component|sram|latches[24][1]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][1]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][1] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][1] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][1] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][1] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][1] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][1] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[15][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[13][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[14][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[12][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[11][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[9][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[10][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[8][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[1][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[2][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[0][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[3][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[21][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[22][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[20][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[23][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[17][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[18][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[16][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[19][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[5][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[6][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[4][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[7][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[31][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[29][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[30][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[28][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[27][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[25][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[26][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][2] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_2),
	.datac(\lpm_ram_dq_component|sram|latches[24][2]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][2] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[15][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[13][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[14][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[12][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[11][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[9][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[10][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[8][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[1][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[2][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[0][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[3][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[21][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[22][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[20][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[23][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[17][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[18][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[16][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[19][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[5][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[6][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[4][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[7][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[31][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[29][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[30][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[28][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[27][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[25][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[26][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][3] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_3),
	.datac(\lpm_ram_dq_component|sram|latches[24][3]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][3]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][3] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[15][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[13][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[14][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[12][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[11][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[9][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[10][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[8][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[1][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[2][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[0][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[3][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[21][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[22][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[20][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[23][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[17][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[18][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[16][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[19][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[5][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[6][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[4][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[7][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[31][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[29][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[30][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[28][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[27][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[25][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[26][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][4] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_4),
	.datac(\lpm_ram_dq_component|sram|latches[24][4]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][4]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][4] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][4] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][4] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][4] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][4] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][4] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[15][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[13][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[14][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[12][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[11][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[9][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[10][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[8][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[1][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[2][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[0][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[3][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[21][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[22][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[20][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[23][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[17][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[18][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[16][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[19][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[5][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[6][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[4][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[7][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[31][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[29][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[30][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[28][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[27][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[25][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[26][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][5] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_5),
	.datac(\lpm_ram_dq_component|sram|latches[24][5]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][5]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][5] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][5] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][5] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][5] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][5] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][5] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[15][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[13][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[14][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[12][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[11][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[9][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[10][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[8][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[1][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[2][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[0][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[3][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[21][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[22][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[20][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[23][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[17][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[18][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[16][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[19][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[5][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[6][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[4][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[7][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[31][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[29][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[30][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[28][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[27][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[25][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[26][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][6] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_6),
	.datac(\lpm_ram_dq_component|sram|latches[24][6]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][6]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][6] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][6] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][6] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][6] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][6] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][6] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[15][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[13][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[14][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[12][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[11][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[9][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[10][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[8][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[1][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[2][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[0][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[3][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[21][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[22][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[20][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[23][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[17][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[18][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[16][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[19][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[5][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[6][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[4][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[7][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[31][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[29][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[30][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[28][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[27][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[25][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[26][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][7] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_7),
	.datac(\lpm_ram_dq_component|sram|latches[24][7]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][7]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][7] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][7] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][7] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][7] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][7] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][7] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[15][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[13][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[14][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[12][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[11][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[9][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[10][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[8][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[1][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[2][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[0][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[3][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[21][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[22][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[20][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[23][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[17][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[18][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[16][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[19][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[5][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[6][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[4][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[7][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[31][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[29][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[30][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[28][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[27][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[25][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[26][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][8] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_8),
	.datac(\lpm_ram_dq_component|sram|latches[24][8]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][8]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][8] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][8] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][8] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][8] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][8] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][8] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[15][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[13][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[14][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[12][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[11][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[9][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[10][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[8][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[1][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[2][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[0][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[3][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[21][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[22][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[20][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[23][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[17][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[18][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[16][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[19][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[5][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[6][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[4][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[7][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[31][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[29][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[30][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[28][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[27][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[25][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[26][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][9] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_9),
	.datac(\lpm_ram_dq_component|sram|latches[24][9]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][9]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][9] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][9] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][9] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][9] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][9] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][9] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[15][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[13][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[14][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[12][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[11][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[9][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[10][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[8][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[1][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[2][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[0][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[3][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[21][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[22][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[20][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[23][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[17][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[18][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[16][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[19][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[5][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[6][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[4][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[7][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[31][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[29][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[30][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[28][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[27][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[25][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[26][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][10] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_10),
	.datac(\lpm_ram_dq_component|sram|latches[24][10]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][10]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][10] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][10] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][10] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][10] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][10] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][10] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[15][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[13][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[14][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[12][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[11][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[9][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[10][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[8][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[1][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[2][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[0][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[3][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[21][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[22][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[20][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[23][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[17][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[18][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[16][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[19][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[5][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[6][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[4][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[7][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[31][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[29][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[30][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[28][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[27][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[25][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[26][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][11] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_11),
	.datac(\lpm_ram_dq_component|sram|latches[24][11]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][11]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][11] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][11] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][11] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][11] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][11] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][11] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[15][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[13][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[14][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[12][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[11][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[9][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[10][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[8][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[1][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[2][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[0][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[3][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[21][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[22][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[20][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[23][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[17][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[18][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[16][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[19][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[5][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[6][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[4][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[7][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[31][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[29][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[30][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[28][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[27][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[25][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[26][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][12] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_12),
	.datac(\lpm_ram_dq_component|sram|latches[24][12]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][12]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][12] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][12] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][12] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][12] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][12] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][12] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[15][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[13][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[14][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[12][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[11][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[9][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[10][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[8][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[1][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[2][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[0][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[3][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[21][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[22][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[20][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[23][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[17][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[18][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[16][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[19][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[5][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[6][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[4][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[7][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[31][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[29][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[30][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[28][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[27][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[25][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[26][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][13] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_13),
	.datac(\lpm_ram_dq_component|sram|latches[24][13]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][13]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][13] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][13] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][13] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][13] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][13] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][13] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[15][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[13][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[14][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[12][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[11][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[9][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[10][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[8][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[1][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[2][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[0][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[3][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[21][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[22][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[20][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[23][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[17][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[18][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[16][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[19][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[5][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[6][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[4][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[7][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[31][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[29][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[30][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[28][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[27][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[25][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[26][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][14] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_14),
	.datac(\lpm_ram_dq_component|sram|latches[24][14]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][14]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][14] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][14] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][14] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][14] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][14] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][14] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[15][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[15][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[15][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[15][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[15][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[15][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[15][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[15][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[15][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[13][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[13][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[13][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[13][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[13][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[13][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[13][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[13][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[13][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[14][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[14][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[14][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[14][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[14][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[14][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[14][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[14][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[14][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[12][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[12][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[12][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[12][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[12][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[12][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[12][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[12][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[12][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[11][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[11][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[11][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[11][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[11][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[11][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[11][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[11][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[11][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[9][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[9][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[9][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[9][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[9][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[9][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[9][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[9][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[9][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[10][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[10][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[10][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[10][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[10][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[10][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[10][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[10][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[10][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[8][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[8][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[8][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[8][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[8][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[8][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[8][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[8][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[8][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[1][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[1][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[1][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[1][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[1][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[1][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[1][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[1][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[1][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[2][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[2][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[2][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[2][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[2][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[2][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[2][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[2][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[2][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[0][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[0][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[0][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[0][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[0][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[0][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[0][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[0][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[0][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[3][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[3][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[3][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[3][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[3][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[3][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[3][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[3][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[3][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[21][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[21][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[21][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[21][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[21][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[21][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[21][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[21][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[21][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[22][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[22][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[22][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[22][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[22][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[22][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[22][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[22][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[22][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[20][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[20][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[20][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[20][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[20][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[20][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[20][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[20][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[20][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[23][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[23][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[23][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[23][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[23][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[23][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[23][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[23][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[23][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[17][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[17][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[17][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[17][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[17][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[17][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[17][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[17][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[17][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[18][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[18][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[18][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[18][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[18][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[18][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[18][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[18][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[18][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[16][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[16][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[16][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[16][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[16][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[16][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[16][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[16][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[16][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[19][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[19][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[19][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[19][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[19][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[19][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[19][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[19][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[19][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[5][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[5][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[5][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[5][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[5][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[5][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[5][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[5][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[5][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[6][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[6][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[6][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[6][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[6][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[6][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[6][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[6][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[6][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[4][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[4][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[4][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[4][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[4][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[4][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[4][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[4][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[4][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[7][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[7][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[7][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[7][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[7][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[7][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[7][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[7][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[7][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[31][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[31][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[31][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[31][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[31][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[31][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[31][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[31][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[31][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[29][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[29][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[29][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[29][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[29][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[29][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[29][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[29][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[29][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[30][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[30][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[30][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[30][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[30][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[30][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[30][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[30][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[30][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[28][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[28][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[28][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[28][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[28][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[28][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[28][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[28][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[28][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[27][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[27][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[27][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[27][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[27][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[27][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[27][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[27][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[27][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[25][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[25][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[25][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[25][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[25][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[25][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[25][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[25][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[25][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[26][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[26][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[26][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[26][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[26][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[26][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[26][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[26][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[26][15] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|latches[24][15] (
	.clk(gnd),
	.dataa(vcc),
	.datab(data_15),
	.datac(\lpm_ram_dq_component|sram|latches[24][15]~combout ),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|latches[24][15]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|latches[24][15] .lut_mask = "ccf0";
defparam \lpm_ram_dq_component|sram|latches[24][15] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|latches[24][15] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|latches[24][15] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|latches[24][15] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|latches[24][15] .synch_mode = "off";

endmodule

module memory_lpm_decode_1 (
	address_0,
	address_1,
	address_2,
	address_4,
	address_3,
	w_anode196w_2,
	w_anode287w_2,
	w_anode165w_3,
	w_anode155w_3,
	w_anode125w_3,
	w_anode114w_3,
	we,
	w_anode135w_3,
	w_anode43w_3,
	w_anode16w_3,
	w_anode226w_3,
	w_anode205w_3,
	w_anode317w_3,
	w_anode185w_3,
	w_anode165w_31,
	w_anode175w_3,
	w_anode155w_31,
	w_anode145w_3,
	w_anode125w_31,
	w_anode114w_31,
	w_anode33w_3,
	w_anode53w_3,
	w_anode256w_3,
	w_anode266w_3,
	w_anode246w_3,
	w_anode276w_3,
	w_anode216w_3,
	w_anode236w_3,
	w_anode73w_3,
	w_anode83w_3,
	w_anode63w_3,
	w_anode93w_3,
	w_anode367w_3,
	w_anode347w_3,
	w_anode357w_3,
	w_anode337w_3,
	w_anode327w_3,
	w_anode307w_3,
	w_anode296w_3)/* synthesis synthesis_greybox=0 */;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_4;
input 	address_3;
output 	w_anode196w_2;
output 	w_anode287w_2;
output 	w_anode165w_3;
output 	w_anode155w_3;
output 	w_anode125w_3;
output 	w_anode114w_3;
input 	we;
output 	w_anode135w_3;
output 	w_anode43w_3;
output 	w_anode16w_3;
output 	w_anode226w_3;
output 	w_anode205w_3;
output 	w_anode317w_3;
output 	w_anode185w_3;
output 	w_anode165w_31;
output 	w_anode175w_3;
output 	w_anode155w_31;
output 	w_anode145w_3;
output 	w_anode125w_31;
output 	w_anode114w_31;
output 	w_anode33w_3;
output 	w_anode53w_3;
output 	w_anode256w_3;
output 	w_anode266w_3;
output 	w_anode246w_3;
output 	w_anode276w_3;
output 	w_anode216w_3;
output 	w_anode236w_3;
output 	w_anode73w_3;
output 	w_anode83w_3;
output 	w_anode63w_3;
output 	w_anode93w_3;
output 	w_anode367w_3;
output 	w_anode347w_3;
output 	w_anode357w_3;
output 	w_anode337w_3;
output 	w_anode327w_3;
output 	w_anode307w_3;
output 	w_anode296w_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



memory_decode_fcf auto_generated(
	.address_0(address_0),
	.address_1(address_1),
	.address_2(address_2),
	.address_4(address_4),
	.address_3(address_3),
	.w_anode196w_2(w_anode196w_2),
	.w_anode287w_2(w_anode287w_2),
	.w_anode165w_3(w_anode165w_3),
	.w_anode155w_3(w_anode155w_3),
	.w_anode125w_3(w_anode125w_3),
	.w_anode114w_3(w_anode114w_3),
	.we(we),
	.w_anode135w_3(w_anode135w_3),
	.w_anode43w_3(w_anode43w_3),
	.w_anode16w_3(w_anode16w_3),
	.w_anode226w_3(w_anode226w_3),
	.w_anode205w_3(w_anode205w_3),
	.w_anode317w_3(w_anode317w_3),
	.w_anode185w_3(w_anode185w_3),
	.w_anode165w_31(w_anode165w_31),
	.w_anode175w_3(w_anode175w_3),
	.w_anode155w_31(w_anode155w_31),
	.w_anode145w_3(w_anode145w_3),
	.w_anode125w_31(w_anode125w_31),
	.w_anode114w_31(w_anode114w_31),
	.w_anode33w_3(w_anode33w_3),
	.w_anode53w_3(w_anode53w_3),
	.w_anode256w_3(w_anode256w_3),
	.w_anode266w_3(w_anode266w_3),
	.w_anode246w_3(w_anode246w_3),
	.w_anode276w_3(w_anode276w_3),
	.w_anode216w_3(w_anode216w_3),
	.w_anode236w_3(w_anode236w_3),
	.w_anode73w_3(w_anode73w_3),
	.w_anode83w_3(w_anode83w_3),
	.w_anode63w_3(w_anode63w_3),
	.w_anode93w_3(w_anode93w_3),
	.w_anode367w_3(w_anode367w_3),
	.w_anode347w_3(w_anode347w_3),
	.w_anode357w_3(w_anode357w_3),
	.w_anode337w_3(w_anode337w_3),
	.w_anode327w_3(w_anode327w_3),
	.w_anode307w_3(w_anode307w_3),
	.w_anode296w_3(w_anode296w_3));

endmodule

module memory_decode_fcf (
	address_0,
	address_1,
	address_2,
	address_4,
	address_3,
	w_anode196w_2,
	w_anode287w_2,
	w_anode165w_3,
	w_anode155w_3,
	w_anode125w_3,
	w_anode114w_3,
	we,
	w_anode135w_3,
	w_anode43w_3,
	w_anode16w_3,
	w_anode226w_3,
	w_anode205w_3,
	w_anode317w_3,
	w_anode185w_3,
	w_anode165w_31,
	w_anode175w_3,
	w_anode155w_31,
	w_anode145w_3,
	w_anode125w_31,
	w_anode114w_31,
	w_anode33w_3,
	w_anode53w_3,
	w_anode256w_3,
	w_anode266w_3,
	w_anode246w_3,
	w_anode276w_3,
	w_anode216w_3,
	w_anode236w_3,
	w_anode73w_3,
	w_anode83w_3,
	w_anode63w_3,
	w_anode93w_3,
	w_anode367w_3,
	w_anode347w_3,
	w_anode357w_3,
	w_anode337w_3,
	w_anode327w_3,
	w_anode307w_3,
	w_anode296w_3)/* synthesis synthesis_greybox=0 */;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_4;
input 	address_3;
output 	w_anode196w_2;
output 	w_anode287w_2;
output 	w_anode165w_3;
output 	w_anode155w_3;
output 	w_anode125w_3;
output 	w_anode114w_3;
input 	we;
output 	w_anode135w_3;
output 	w_anode43w_3;
output 	w_anode16w_3;
output 	w_anode226w_3;
output 	w_anode205w_3;
output 	w_anode317w_3;
output 	w_anode185w_3;
output 	w_anode165w_31;
output 	w_anode175w_3;
output 	w_anode155w_31;
output 	w_anode145w_3;
output 	w_anode125w_31;
output 	w_anode114w_31;
output 	w_anode33w_3;
output 	w_anode53w_3;
output 	w_anode256w_3;
output 	w_anode266w_3;
output 	w_anode246w_3;
output 	w_anode276w_3;
output 	w_anode216w_3;
output 	w_anode236w_3;
output 	w_anode73w_3;
output 	w_anode83w_3;
output 	w_anode63w_3;
output 	w_anode93w_3;
output 	w_anode367w_3;
output 	w_anode347w_3;
output 	w_anode357w_3;
output 	w_anode337w_3;
output 	w_anode327w_3;
output 	w_anode307w_3;
output 	w_anode296w_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ;
wire \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ;


maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 (
	.clk(gnd),
	.dataa(address_4),
	.datab(vcc),
	.datac(vcc),
	.datad(address_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode196w_2),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 .lut_mask = "00aa";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~0 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_4),
	.datac(vcc),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode287w_2),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 .lut_mask = "8888";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~0 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(vcc),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode165w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 .lut_mask = "8888";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3]~2 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 (
	.clk(gnd),
	.dataa(address_2),
	.datab(vcc),
	.datac(vcc),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode155w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 .lut_mask = "00aa";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3]~2 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 (
	.clk(gnd),
	.dataa(address_0),
	.datab(vcc),
	.datac(vcc),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode125w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 .lut_mask = "00aa";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3]~2 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 (
	.clk(gnd),
	.dataa(vcc),
	.datab(vcc),
	.datac(address_0),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode114w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 .lut_mask = "000f";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3]~2 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] (
	.clk(gnd),
	.dataa(address_1),
	.datab(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.datac(address_0),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode135w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] .lut_mask = "0008";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode135w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] (
	.clk(gnd),
	.dataa(address_1),
	.datab(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.datac(address_0),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode43w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] .lut_mask = "0008";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode43w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.datab(address_0),
	.datac(address_1),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode16w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] .lut_mask = "0002";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode16w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] (
	.clk(gnd),
	.dataa(address_1),
	.datab(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.datac(address_0),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode226w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] .lut_mask = "0008";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode226w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.datab(address_0),
	.datac(address_1),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode205w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] .lut_mask = "0002";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode205w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] (
	.clk(gnd),
	.dataa(address_1),
	.datab(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.datac(address_0),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode317w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] .lut_mask = "0008";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode317w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode185w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] .lut_mask = "8000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode185w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode165w_31),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] .lut_mask = "0080";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode165w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode175w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode175w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode155w_31),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode155w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode145w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode145w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode125w_31),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode125w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode114w_31),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] .lut_mask = "0010";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode114w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode33w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode33w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode53w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode53w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode256w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] .lut_mask = "0080";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode256w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode266w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode266w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode246w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode246w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode276w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] .lut_mask = "8000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode276w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode216w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode216w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode236w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode236w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode73w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] .lut_mask = "0080";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode73w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode83w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode83w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode63w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode63w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode93w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] .lut_mask = "8000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode93w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode367w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] .lut_mask = "8000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode367w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode347w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] .lut_mask = "0080";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode347w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode357w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode357w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] (
	.clk(gnd),
	.dataa(address_2),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode337w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode337w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(address_1),
	.datad(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode327w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] .lut_mask = "2000";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode327w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode307w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] .lut_mask = "0020";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode307w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] (
	.clk(gnd),
	.dataa(address_0),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(w_anode296w_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] .lut_mask = "0010";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode296w[3] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] (
	.clk(gnd),
	.dataa(address_3),
	.datab(we),
	.datac(vcc),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] .lut_mask = "0088";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode105w[2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] (
	.clk(gnd),
	.dataa(we),
	.datab(vcc),
	.datac(address_3),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] .lut_mask = "000a";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode3w[2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] (
	.clk(gnd),
	.dataa(address_4),
	.datab(we),
	.datac(vcc),
	.datad(address_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] .lut_mask = "0088";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode196w[2] .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_4),
	.datac(we),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2]~combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] .lut_mask = "8080";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|decode|auto_generated|w_anode287w[2] .synch_mode = "off";

endmodule

module memory_lpm_mux_1 (
	address_0,
	address_1,
	address_2,
	address_4,
	address_3,
	w_anode196w_2,
	w_anode287w_2,
	w_anode165w_3,
	w_anode155w_3,
	w_anode125w_3,
	w_anode114w_3,
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	latches_0_15,
	latches_0_13,
	latches_0_14,
	latches_0_12,
	latches_0_11,
	latches_0_9,
	latches_0_10,
	latches_0_8,
	latches_0_1,
	latches_0_2,
	latches_0_0,
	latches_0_3,
	latches_0_21,
	latches_0_22,
	latches_0_20,
	latches_0_23,
	latches_0_17,
	latches_0_18,
	latches_0_16,
	latches_0_19,
	latches_0_5,
	latches_0_6,
	latches_0_4,
	latches_0_7,
	latches_0_31,
	latches_0_29,
	latches_0_30,
	latches_0_28,
	latches_0_27,
	latches_0_25,
	latches_0_26,
	latches_0_24,
	latches_1_15,
	latches_1_13,
	latches_1_14,
	latches_1_12,
	latches_1_11,
	latches_1_9,
	latches_1_10,
	latches_1_8,
	latches_1_1,
	latches_1_2,
	latches_1_0,
	latches_1_3,
	latches_1_21,
	latches_1_22,
	latches_1_20,
	latches_1_23,
	latches_1_17,
	latches_1_18,
	latches_1_16,
	latches_1_19,
	latches_1_5,
	latches_1_6,
	latches_1_4,
	latches_1_7,
	latches_1_31,
	latches_1_29,
	latches_1_30,
	latches_1_28,
	latches_1_27,
	latches_1_25,
	latches_1_26,
	latches_1_24,
	latches_2_15,
	latches_2_13,
	latches_2_14,
	latches_2_12,
	latches_2_11,
	latches_2_9,
	latches_2_10,
	latches_2_8,
	latches_2_1,
	latches_2_2,
	latches_2_0,
	latches_2_3,
	latches_2_21,
	latches_2_22,
	latches_2_20,
	latches_2_23,
	latches_2_17,
	latches_2_18,
	latches_2_16,
	latches_2_19,
	latches_2_5,
	latches_2_6,
	latches_2_4,
	latches_2_7,
	latches_2_31,
	latches_2_29,
	latches_2_30,
	latches_2_28,
	latches_2_27,
	latches_2_25,
	latches_2_26,
	latches_2_24,
	latches_3_15,
	latches_3_13,
	latches_3_14,
	latches_3_12,
	latches_3_11,
	latches_3_9,
	latches_3_10,
	latches_3_8,
	latches_3_1,
	latches_3_2,
	latches_3_0,
	latches_3_3,
	latches_3_21,
	latches_3_22,
	latches_3_20,
	latches_3_23,
	latches_3_17,
	latches_3_18,
	latches_3_16,
	latches_3_19,
	latches_3_5,
	latches_3_6,
	latches_3_4,
	latches_3_7,
	latches_3_31,
	latches_3_29,
	latches_3_30,
	latches_3_28,
	latches_3_27,
	latches_3_25,
	latches_3_26,
	latches_3_24,
	latches_4_15,
	latches_4_13,
	latches_4_14,
	latches_4_12,
	latches_4_11,
	latches_4_9,
	latches_4_10,
	latches_4_8,
	latches_4_1,
	latches_4_2,
	latches_4_0,
	latches_4_3,
	latches_4_21,
	latches_4_22,
	latches_4_20,
	latches_4_23,
	latches_4_17,
	latches_4_18,
	latches_4_16,
	latches_4_19,
	latches_4_5,
	latches_4_6,
	latches_4_4,
	latches_4_7,
	latches_4_31,
	latches_4_29,
	latches_4_30,
	latches_4_28,
	latches_4_27,
	latches_4_25,
	latches_4_26,
	latches_4_24,
	latches_5_15,
	latches_5_13,
	latches_5_14,
	latches_5_12,
	latches_5_11,
	latches_5_9,
	latches_5_10,
	latches_5_8,
	latches_5_1,
	latches_5_2,
	latches_5_0,
	latches_5_3,
	latches_5_21,
	latches_5_22,
	latches_5_20,
	latches_5_23,
	latches_5_17,
	latches_5_18,
	latches_5_16,
	latches_5_19,
	latches_5_5,
	latches_5_6,
	latches_5_4,
	latches_5_7,
	latches_5_31,
	latches_5_29,
	latches_5_30,
	latches_5_28,
	latches_5_27,
	latches_5_25,
	latches_5_26,
	latches_5_24,
	latches_6_15,
	latches_6_13,
	latches_6_14,
	latches_6_12,
	latches_6_11,
	latches_6_9,
	latches_6_10,
	latches_6_8,
	latches_6_1,
	latches_6_2,
	latches_6_0,
	latches_6_3,
	latches_6_21,
	latches_6_22,
	latches_6_20,
	latches_6_23,
	latches_6_17,
	latches_6_18,
	latches_6_16,
	latches_6_19,
	latches_6_5,
	latches_6_6,
	latches_6_4,
	latches_6_7,
	latches_6_31,
	latches_6_29,
	latches_6_30,
	latches_6_28,
	latches_6_27,
	latches_6_25,
	latches_6_26,
	latches_6_24,
	latches_7_15,
	latches_7_13,
	latches_7_14,
	latches_7_12,
	latches_7_11,
	latches_7_9,
	latches_7_10,
	latches_7_8,
	latches_7_1,
	latches_7_2,
	latches_7_0,
	latches_7_3,
	latches_7_21,
	latches_7_22,
	latches_7_20,
	latches_7_23,
	latches_7_17,
	latches_7_18,
	latches_7_16,
	latches_7_19,
	latches_7_5,
	latches_7_6,
	latches_7_4,
	latches_7_7,
	latches_7_31,
	latches_7_29,
	latches_7_30,
	latches_7_28,
	latches_7_27,
	latches_7_25,
	latches_7_26,
	latches_7_24,
	latches_8_15,
	latches_8_13,
	latches_8_14,
	latches_8_12,
	latches_8_11,
	latches_8_9,
	latches_8_10,
	latches_8_8,
	latches_8_1,
	latches_8_2,
	latches_8_0,
	latches_8_3,
	latches_8_21,
	latches_8_22,
	latches_8_20,
	latches_8_23,
	latches_8_17,
	latches_8_18,
	latches_8_16,
	latches_8_19,
	latches_8_5,
	latches_8_6,
	latches_8_4,
	latches_8_7,
	latches_8_31,
	latches_8_29,
	latches_8_30,
	latches_8_28,
	latches_8_27,
	latches_8_25,
	latches_8_26,
	latches_8_24,
	latches_9_15,
	latches_9_13,
	latches_9_14,
	latches_9_12,
	latches_9_11,
	latches_9_9,
	latches_9_10,
	latches_9_8,
	latches_9_1,
	latches_9_2,
	latches_9_0,
	latches_9_3,
	latches_9_21,
	latches_9_22,
	latches_9_20,
	latches_9_23,
	latches_9_17,
	latches_9_18,
	latches_9_16,
	latches_9_19,
	latches_9_5,
	latches_9_6,
	latches_9_4,
	latches_9_7,
	latches_9_31,
	latches_9_29,
	latches_9_30,
	latches_9_28,
	latches_9_27,
	latches_9_25,
	latches_9_26,
	latches_9_24,
	latches_10_15,
	latches_10_13,
	latches_10_14,
	latches_10_12,
	latches_10_11,
	latches_10_9,
	latches_10_10,
	latches_10_8,
	latches_10_1,
	latches_10_2,
	latches_10_0,
	latches_10_3,
	latches_10_21,
	latches_10_22,
	latches_10_20,
	latches_10_23,
	latches_10_17,
	latches_10_18,
	latches_10_16,
	latches_10_19,
	latches_10_5,
	latches_10_6,
	latches_10_4,
	latches_10_7,
	latches_10_31,
	latches_10_29,
	latches_10_30,
	latches_10_28,
	latches_10_27,
	latches_10_25,
	latches_10_26,
	latches_10_24,
	latches_11_15,
	latches_11_13,
	latches_11_14,
	latches_11_12,
	latches_11_11,
	latches_11_9,
	latches_11_10,
	latches_11_8,
	latches_11_1,
	latches_11_2,
	latches_11_0,
	latches_11_3,
	latches_11_21,
	latches_11_22,
	latches_11_20,
	latches_11_23,
	latches_11_17,
	latches_11_18,
	latches_11_16,
	latches_11_19,
	latches_11_5,
	latches_11_6,
	latches_11_4,
	latches_11_7,
	latches_11_31,
	latches_11_29,
	latches_11_30,
	latches_11_28,
	latches_11_27,
	latches_11_25,
	latches_11_26,
	latches_11_24,
	latches_12_15,
	latches_12_13,
	latches_12_14,
	latches_12_12,
	latches_12_11,
	latches_12_9,
	latches_12_10,
	latches_12_8,
	latches_12_1,
	latches_12_2,
	latches_12_0,
	latches_12_3,
	latches_12_21,
	latches_12_22,
	latches_12_20,
	latches_12_23,
	latches_12_17,
	latches_12_18,
	latches_12_16,
	latches_12_19,
	latches_12_5,
	latches_12_6,
	latches_12_4,
	latches_12_7,
	latches_12_31,
	latches_12_29,
	latches_12_30,
	latches_12_28,
	latches_12_27,
	latches_12_25,
	latches_12_26,
	latches_12_24,
	latches_13_15,
	latches_13_13,
	latches_13_14,
	latches_13_12,
	latches_13_11,
	latches_13_9,
	latches_13_10,
	latches_13_8,
	latches_13_1,
	latches_13_2,
	latches_13_0,
	latches_13_3,
	latches_13_21,
	latches_13_22,
	latches_13_20,
	latches_13_23,
	latches_13_17,
	latches_13_18,
	latches_13_16,
	latches_13_19,
	latches_13_5,
	latches_13_6,
	latches_13_4,
	latches_13_7,
	latches_13_31,
	latches_13_29,
	latches_13_30,
	latches_13_28,
	latches_13_27,
	latches_13_25,
	latches_13_26,
	latches_13_24,
	latches_14_15,
	latches_14_13,
	latches_14_14,
	latches_14_12,
	latches_14_11,
	latches_14_9,
	latches_14_10,
	latches_14_8,
	latches_14_1,
	latches_14_2,
	latches_14_0,
	latches_14_3,
	latches_14_21,
	latches_14_22,
	latches_14_20,
	latches_14_23,
	latches_14_17,
	latches_14_18,
	latches_14_16,
	latches_14_19,
	latches_14_5,
	latches_14_6,
	latches_14_4,
	latches_14_7,
	latches_14_31,
	latches_14_29,
	latches_14_30,
	latches_14_28,
	latches_14_27,
	latches_14_25,
	latches_14_26,
	latches_14_24,
	latches_15_15,
	latches_15_13,
	latches_15_14,
	latches_15_12,
	latches_15_11,
	latches_15_9,
	latches_15_10,
	latches_15_8,
	latches_15_1,
	latches_15_2,
	latches_15_0,
	latches_15_3,
	latches_15_21,
	latches_15_22,
	latches_15_20,
	latches_15_23,
	latches_15_17,
	latches_15_18,
	latches_15_16,
	latches_15_19,
	latches_15_5,
	latches_15_6,
	latches_15_4,
	latches_15_7,
	latches_15_31,
	latches_15_29,
	latches_15_30,
	latches_15_28,
	latches_15_27,
	latches_15_25,
	latches_15_26,
	latches_15_24)/* synthesis synthesis_greybox=0 */;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_4;
input 	address_3;
input 	w_anode196w_2;
input 	w_anode287w_2;
input 	w_anode165w_3;
input 	w_anode155w_3;
input 	w_anode125w_3;
input 	w_anode114w_3;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
input 	latches_0_15;
input 	latches_0_13;
input 	latches_0_14;
input 	latches_0_12;
input 	latches_0_11;
input 	latches_0_9;
input 	latches_0_10;
input 	latches_0_8;
input 	latches_0_1;
input 	latches_0_2;
input 	latches_0_0;
input 	latches_0_3;
input 	latches_0_21;
input 	latches_0_22;
input 	latches_0_20;
input 	latches_0_23;
input 	latches_0_17;
input 	latches_0_18;
input 	latches_0_16;
input 	latches_0_19;
input 	latches_0_5;
input 	latches_0_6;
input 	latches_0_4;
input 	latches_0_7;
input 	latches_0_31;
input 	latches_0_29;
input 	latches_0_30;
input 	latches_0_28;
input 	latches_0_27;
input 	latches_0_25;
input 	latches_0_26;
input 	latches_0_24;
input 	latches_1_15;
input 	latches_1_13;
input 	latches_1_14;
input 	latches_1_12;
input 	latches_1_11;
input 	latches_1_9;
input 	latches_1_10;
input 	latches_1_8;
input 	latches_1_1;
input 	latches_1_2;
input 	latches_1_0;
input 	latches_1_3;
input 	latches_1_21;
input 	latches_1_22;
input 	latches_1_20;
input 	latches_1_23;
input 	latches_1_17;
input 	latches_1_18;
input 	latches_1_16;
input 	latches_1_19;
input 	latches_1_5;
input 	latches_1_6;
input 	latches_1_4;
input 	latches_1_7;
input 	latches_1_31;
input 	latches_1_29;
input 	latches_1_30;
input 	latches_1_28;
input 	latches_1_27;
input 	latches_1_25;
input 	latches_1_26;
input 	latches_1_24;
input 	latches_2_15;
input 	latches_2_13;
input 	latches_2_14;
input 	latches_2_12;
input 	latches_2_11;
input 	latches_2_9;
input 	latches_2_10;
input 	latches_2_8;
input 	latches_2_1;
input 	latches_2_2;
input 	latches_2_0;
input 	latches_2_3;
input 	latches_2_21;
input 	latches_2_22;
input 	latches_2_20;
input 	latches_2_23;
input 	latches_2_17;
input 	latches_2_18;
input 	latches_2_16;
input 	latches_2_19;
input 	latches_2_5;
input 	latches_2_6;
input 	latches_2_4;
input 	latches_2_7;
input 	latches_2_31;
input 	latches_2_29;
input 	latches_2_30;
input 	latches_2_28;
input 	latches_2_27;
input 	latches_2_25;
input 	latches_2_26;
input 	latches_2_24;
input 	latches_3_15;
input 	latches_3_13;
input 	latches_3_14;
input 	latches_3_12;
input 	latches_3_11;
input 	latches_3_9;
input 	latches_3_10;
input 	latches_3_8;
input 	latches_3_1;
input 	latches_3_2;
input 	latches_3_0;
input 	latches_3_3;
input 	latches_3_21;
input 	latches_3_22;
input 	latches_3_20;
input 	latches_3_23;
input 	latches_3_17;
input 	latches_3_18;
input 	latches_3_16;
input 	latches_3_19;
input 	latches_3_5;
input 	latches_3_6;
input 	latches_3_4;
input 	latches_3_7;
input 	latches_3_31;
input 	latches_3_29;
input 	latches_3_30;
input 	latches_3_28;
input 	latches_3_27;
input 	latches_3_25;
input 	latches_3_26;
input 	latches_3_24;
input 	latches_4_15;
input 	latches_4_13;
input 	latches_4_14;
input 	latches_4_12;
input 	latches_4_11;
input 	latches_4_9;
input 	latches_4_10;
input 	latches_4_8;
input 	latches_4_1;
input 	latches_4_2;
input 	latches_4_0;
input 	latches_4_3;
input 	latches_4_21;
input 	latches_4_22;
input 	latches_4_20;
input 	latches_4_23;
input 	latches_4_17;
input 	latches_4_18;
input 	latches_4_16;
input 	latches_4_19;
input 	latches_4_5;
input 	latches_4_6;
input 	latches_4_4;
input 	latches_4_7;
input 	latches_4_31;
input 	latches_4_29;
input 	latches_4_30;
input 	latches_4_28;
input 	latches_4_27;
input 	latches_4_25;
input 	latches_4_26;
input 	latches_4_24;
input 	latches_5_15;
input 	latches_5_13;
input 	latches_5_14;
input 	latches_5_12;
input 	latches_5_11;
input 	latches_5_9;
input 	latches_5_10;
input 	latches_5_8;
input 	latches_5_1;
input 	latches_5_2;
input 	latches_5_0;
input 	latches_5_3;
input 	latches_5_21;
input 	latches_5_22;
input 	latches_5_20;
input 	latches_5_23;
input 	latches_5_17;
input 	latches_5_18;
input 	latches_5_16;
input 	latches_5_19;
input 	latches_5_5;
input 	latches_5_6;
input 	latches_5_4;
input 	latches_5_7;
input 	latches_5_31;
input 	latches_5_29;
input 	latches_5_30;
input 	latches_5_28;
input 	latches_5_27;
input 	latches_5_25;
input 	latches_5_26;
input 	latches_5_24;
input 	latches_6_15;
input 	latches_6_13;
input 	latches_6_14;
input 	latches_6_12;
input 	latches_6_11;
input 	latches_6_9;
input 	latches_6_10;
input 	latches_6_8;
input 	latches_6_1;
input 	latches_6_2;
input 	latches_6_0;
input 	latches_6_3;
input 	latches_6_21;
input 	latches_6_22;
input 	latches_6_20;
input 	latches_6_23;
input 	latches_6_17;
input 	latches_6_18;
input 	latches_6_16;
input 	latches_6_19;
input 	latches_6_5;
input 	latches_6_6;
input 	latches_6_4;
input 	latches_6_7;
input 	latches_6_31;
input 	latches_6_29;
input 	latches_6_30;
input 	latches_6_28;
input 	latches_6_27;
input 	latches_6_25;
input 	latches_6_26;
input 	latches_6_24;
input 	latches_7_15;
input 	latches_7_13;
input 	latches_7_14;
input 	latches_7_12;
input 	latches_7_11;
input 	latches_7_9;
input 	latches_7_10;
input 	latches_7_8;
input 	latches_7_1;
input 	latches_7_2;
input 	latches_7_0;
input 	latches_7_3;
input 	latches_7_21;
input 	latches_7_22;
input 	latches_7_20;
input 	latches_7_23;
input 	latches_7_17;
input 	latches_7_18;
input 	latches_7_16;
input 	latches_7_19;
input 	latches_7_5;
input 	latches_7_6;
input 	latches_7_4;
input 	latches_7_7;
input 	latches_7_31;
input 	latches_7_29;
input 	latches_7_30;
input 	latches_7_28;
input 	latches_7_27;
input 	latches_7_25;
input 	latches_7_26;
input 	latches_7_24;
input 	latches_8_15;
input 	latches_8_13;
input 	latches_8_14;
input 	latches_8_12;
input 	latches_8_11;
input 	latches_8_9;
input 	latches_8_10;
input 	latches_8_8;
input 	latches_8_1;
input 	latches_8_2;
input 	latches_8_0;
input 	latches_8_3;
input 	latches_8_21;
input 	latches_8_22;
input 	latches_8_20;
input 	latches_8_23;
input 	latches_8_17;
input 	latches_8_18;
input 	latches_8_16;
input 	latches_8_19;
input 	latches_8_5;
input 	latches_8_6;
input 	latches_8_4;
input 	latches_8_7;
input 	latches_8_31;
input 	latches_8_29;
input 	latches_8_30;
input 	latches_8_28;
input 	latches_8_27;
input 	latches_8_25;
input 	latches_8_26;
input 	latches_8_24;
input 	latches_9_15;
input 	latches_9_13;
input 	latches_9_14;
input 	latches_9_12;
input 	latches_9_11;
input 	latches_9_9;
input 	latches_9_10;
input 	latches_9_8;
input 	latches_9_1;
input 	latches_9_2;
input 	latches_9_0;
input 	latches_9_3;
input 	latches_9_21;
input 	latches_9_22;
input 	latches_9_20;
input 	latches_9_23;
input 	latches_9_17;
input 	latches_9_18;
input 	latches_9_16;
input 	latches_9_19;
input 	latches_9_5;
input 	latches_9_6;
input 	latches_9_4;
input 	latches_9_7;
input 	latches_9_31;
input 	latches_9_29;
input 	latches_9_30;
input 	latches_9_28;
input 	latches_9_27;
input 	latches_9_25;
input 	latches_9_26;
input 	latches_9_24;
input 	latches_10_15;
input 	latches_10_13;
input 	latches_10_14;
input 	latches_10_12;
input 	latches_10_11;
input 	latches_10_9;
input 	latches_10_10;
input 	latches_10_8;
input 	latches_10_1;
input 	latches_10_2;
input 	latches_10_0;
input 	latches_10_3;
input 	latches_10_21;
input 	latches_10_22;
input 	latches_10_20;
input 	latches_10_23;
input 	latches_10_17;
input 	latches_10_18;
input 	latches_10_16;
input 	latches_10_19;
input 	latches_10_5;
input 	latches_10_6;
input 	latches_10_4;
input 	latches_10_7;
input 	latches_10_31;
input 	latches_10_29;
input 	latches_10_30;
input 	latches_10_28;
input 	latches_10_27;
input 	latches_10_25;
input 	latches_10_26;
input 	latches_10_24;
input 	latches_11_15;
input 	latches_11_13;
input 	latches_11_14;
input 	latches_11_12;
input 	latches_11_11;
input 	latches_11_9;
input 	latches_11_10;
input 	latches_11_8;
input 	latches_11_1;
input 	latches_11_2;
input 	latches_11_0;
input 	latches_11_3;
input 	latches_11_21;
input 	latches_11_22;
input 	latches_11_20;
input 	latches_11_23;
input 	latches_11_17;
input 	latches_11_18;
input 	latches_11_16;
input 	latches_11_19;
input 	latches_11_5;
input 	latches_11_6;
input 	latches_11_4;
input 	latches_11_7;
input 	latches_11_31;
input 	latches_11_29;
input 	latches_11_30;
input 	latches_11_28;
input 	latches_11_27;
input 	latches_11_25;
input 	latches_11_26;
input 	latches_11_24;
input 	latches_12_15;
input 	latches_12_13;
input 	latches_12_14;
input 	latches_12_12;
input 	latches_12_11;
input 	latches_12_9;
input 	latches_12_10;
input 	latches_12_8;
input 	latches_12_1;
input 	latches_12_2;
input 	latches_12_0;
input 	latches_12_3;
input 	latches_12_21;
input 	latches_12_22;
input 	latches_12_20;
input 	latches_12_23;
input 	latches_12_17;
input 	latches_12_18;
input 	latches_12_16;
input 	latches_12_19;
input 	latches_12_5;
input 	latches_12_6;
input 	latches_12_4;
input 	latches_12_7;
input 	latches_12_31;
input 	latches_12_29;
input 	latches_12_30;
input 	latches_12_28;
input 	latches_12_27;
input 	latches_12_25;
input 	latches_12_26;
input 	latches_12_24;
input 	latches_13_15;
input 	latches_13_13;
input 	latches_13_14;
input 	latches_13_12;
input 	latches_13_11;
input 	latches_13_9;
input 	latches_13_10;
input 	latches_13_8;
input 	latches_13_1;
input 	latches_13_2;
input 	latches_13_0;
input 	latches_13_3;
input 	latches_13_21;
input 	latches_13_22;
input 	latches_13_20;
input 	latches_13_23;
input 	latches_13_17;
input 	latches_13_18;
input 	latches_13_16;
input 	latches_13_19;
input 	latches_13_5;
input 	latches_13_6;
input 	latches_13_4;
input 	latches_13_7;
input 	latches_13_31;
input 	latches_13_29;
input 	latches_13_30;
input 	latches_13_28;
input 	latches_13_27;
input 	latches_13_25;
input 	latches_13_26;
input 	latches_13_24;
input 	latches_14_15;
input 	latches_14_13;
input 	latches_14_14;
input 	latches_14_12;
input 	latches_14_11;
input 	latches_14_9;
input 	latches_14_10;
input 	latches_14_8;
input 	latches_14_1;
input 	latches_14_2;
input 	latches_14_0;
input 	latches_14_3;
input 	latches_14_21;
input 	latches_14_22;
input 	latches_14_20;
input 	latches_14_23;
input 	latches_14_17;
input 	latches_14_18;
input 	latches_14_16;
input 	latches_14_19;
input 	latches_14_5;
input 	latches_14_6;
input 	latches_14_4;
input 	latches_14_7;
input 	latches_14_31;
input 	latches_14_29;
input 	latches_14_30;
input 	latches_14_28;
input 	latches_14_27;
input 	latches_14_25;
input 	latches_14_26;
input 	latches_14_24;
input 	latches_15_15;
input 	latches_15_13;
input 	latches_15_14;
input 	latches_15_12;
input 	latches_15_11;
input 	latches_15_9;
input 	latches_15_10;
input 	latches_15_8;
input 	latches_15_1;
input 	latches_15_2;
input 	latches_15_0;
input 	latches_15_3;
input 	latches_15_21;
input 	latches_15_22;
input 	latches_15_20;
input 	latches_15_23;
input 	latches_15_17;
input 	latches_15_18;
input 	latches_15_16;
input 	latches_15_19;
input 	latches_15_5;
input 	latches_15_6;
input 	latches_15_4;
input 	latches_15_7;
input 	latches_15_31;
input 	latches_15_29;
input 	latches_15_30;
input 	latches_15_28;
input 	latches_15_27;
input 	latches_15_25;
input 	latches_15_26;
input 	latches_15_24;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



memory_mux_v9c auto_generated(
	.address_0(address_0),
	.address_1(address_1),
	.address_2(address_2),
	.address_4(address_4),
	.address_3(address_3),
	.w_anode196w_2(w_anode196w_2),
	.w_anode287w_2(w_anode287w_2),
	.w_anode165w_3(w_anode165w_3),
	.w_anode155w_3(w_anode155w_3),
	.w_anode125w_3(w_anode125w_3),
	.w_anode114w_3(w_anode114w_3),
	.result_node_0(result_node_0),
	.result_node_1(result_node_1),
	.result_node_2(result_node_2),
	.result_node_3(result_node_3),
	.result_node_4(result_node_4),
	.result_node_5(result_node_5),
	.result_node_6(result_node_6),
	.result_node_7(result_node_7),
	.result_node_8(result_node_8),
	.result_node_9(result_node_9),
	.result_node_10(result_node_10),
	.result_node_11(result_node_11),
	.result_node_12(result_node_12),
	.result_node_13(result_node_13),
	.result_node_14(result_node_14),
	.result_node_15(result_node_15),
	.latches_0_15(latches_0_15),
	.latches_0_13(latches_0_13),
	.latches_0_14(latches_0_14),
	.latches_0_12(latches_0_12),
	.latches_0_11(latches_0_11),
	.latches_0_9(latches_0_9),
	.latches_0_10(latches_0_10),
	.latches_0_8(latches_0_8),
	.latches_0_1(latches_0_1),
	.latches_0_2(latches_0_2),
	.latches_0_0(latches_0_0),
	.latches_0_3(latches_0_3),
	.latches_0_21(latches_0_21),
	.latches_0_22(latches_0_22),
	.latches_0_20(latches_0_20),
	.latches_0_23(latches_0_23),
	.latches_0_17(latches_0_17),
	.latches_0_18(latches_0_18),
	.latches_0_16(latches_0_16),
	.latches_0_19(latches_0_19),
	.latches_0_5(latches_0_5),
	.latches_0_6(latches_0_6),
	.latches_0_4(latches_0_4),
	.latches_0_7(latches_0_7),
	.latches_0_31(latches_0_31),
	.latches_0_29(latches_0_29),
	.latches_0_30(latches_0_30),
	.latches_0_28(latches_0_28),
	.latches_0_27(latches_0_27),
	.latches_0_25(latches_0_25),
	.latches_0_26(latches_0_26),
	.latches_0_24(latches_0_24),
	.latches_1_15(latches_1_15),
	.latches_1_13(latches_1_13),
	.latches_1_14(latches_1_14),
	.latches_1_12(latches_1_12),
	.latches_1_11(latches_1_11),
	.latches_1_9(latches_1_9),
	.latches_1_10(latches_1_10),
	.latches_1_8(latches_1_8),
	.latches_1_1(latches_1_1),
	.latches_1_2(latches_1_2),
	.latches_1_0(latches_1_0),
	.latches_1_3(latches_1_3),
	.latches_1_21(latches_1_21),
	.latches_1_22(latches_1_22),
	.latches_1_20(latches_1_20),
	.latches_1_23(latches_1_23),
	.latches_1_17(latches_1_17),
	.latches_1_18(latches_1_18),
	.latches_1_16(latches_1_16),
	.latches_1_19(latches_1_19),
	.latches_1_5(latches_1_5),
	.latches_1_6(latches_1_6),
	.latches_1_4(latches_1_4),
	.latches_1_7(latches_1_7),
	.latches_1_31(latches_1_31),
	.latches_1_29(latches_1_29),
	.latches_1_30(latches_1_30),
	.latches_1_28(latches_1_28),
	.latches_1_27(latches_1_27),
	.latches_1_25(latches_1_25),
	.latches_1_26(latches_1_26),
	.latches_1_24(latches_1_24),
	.latches_2_15(latches_2_15),
	.latches_2_13(latches_2_13),
	.latches_2_14(latches_2_14),
	.latches_2_12(latches_2_12),
	.latches_2_11(latches_2_11),
	.latches_2_9(latches_2_9),
	.latches_2_10(latches_2_10),
	.latches_2_8(latches_2_8),
	.latches_2_1(latches_2_1),
	.latches_2_2(latches_2_2),
	.latches_2_0(latches_2_0),
	.latches_2_3(latches_2_3),
	.latches_2_21(latches_2_21),
	.latches_2_22(latches_2_22),
	.latches_2_20(latches_2_20),
	.latches_2_23(latches_2_23),
	.latches_2_17(latches_2_17),
	.latches_2_18(latches_2_18),
	.latches_2_16(latches_2_16),
	.latches_2_19(latches_2_19),
	.latches_2_5(latches_2_5),
	.latches_2_6(latches_2_6),
	.latches_2_4(latches_2_4),
	.latches_2_7(latches_2_7),
	.latches_2_31(latches_2_31),
	.latches_2_29(latches_2_29),
	.latches_2_30(latches_2_30),
	.latches_2_28(latches_2_28),
	.latches_2_27(latches_2_27),
	.latches_2_25(latches_2_25),
	.latches_2_26(latches_2_26),
	.latches_2_24(latches_2_24),
	.latches_3_15(latches_3_15),
	.latches_3_13(latches_3_13),
	.latches_3_14(latches_3_14),
	.latches_3_12(latches_3_12),
	.latches_3_11(latches_3_11),
	.latches_3_9(latches_3_9),
	.latches_3_10(latches_3_10),
	.latches_3_8(latches_3_8),
	.latches_3_1(latches_3_1),
	.latches_3_2(latches_3_2),
	.latches_3_0(latches_3_0),
	.latches_3_3(latches_3_3),
	.latches_3_21(latches_3_21),
	.latches_3_22(latches_3_22),
	.latches_3_20(latches_3_20),
	.latches_3_23(latches_3_23),
	.latches_3_17(latches_3_17),
	.latches_3_18(latches_3_18),
	.latches_3_16(latches_3_16),
	.latches_3_19(latches_3_19),
	.latches_3_5(latches_3_5),
	.latches_3_6(latches_3_6),
	.latches_3_4(latches_3_4),
	.latches_3_7(latches_3_7),
	.latches_3_31(latches_3_31),
	.latches_3_29(latches_3_29),
	.latches_3_30(latches_3_30),
	.latches_3_28(latches_3_28),
	.latches_3_27(latches_3_27),
	.latches_3_25(latches_3_25),
	.latches_3_26(latches_3_26),
	.latches_3_24(latches_3_24),
	.latches_4_15(latches_4_15),
	.latches_4_13(latches_4_13),
	.latches_4_14(latches_4_14),
	.latches_4_12(latches_4_12),
	.latches_4_11(latches_4_11),
	.latches_4_9(latches_4_9),
	.latches_4_10(latches_4_10),
	.latches_4_8(latches_4_8),
	.latches_4_1(latches_4_1),
	.latches_4_2(latches_4_2),
	.latches_4_0(latches_4_0),
	.latches_4_3(latches_4_3),
	.latches_4_21(latches_4_21),
	.latches_4_22(latches_4_22),
	.latches_4_20(latches_4_20),
	.latches_4_23(latches_4_23),
	.latches_4_17(latches_4_17),
	.latches_4_18(latches_4_18),
	.latches_4_16(latches_4_16),
	.latches_4_19(latches_4_19),
	.latches_4_5(latches_4_5),
	.latches_4_6(latches_4_6),
	.latches_4_4(latches_4_4),
	.latches_4_7(latches_4_7),
	.latches_4_31(latches_4_31),
	.latches_4_29(latches_4_29),
	.latches_4_30(latches_4_30),
	.latches_4_28(latches_4_28),
	.latches_4_27(latches_4_27),
	.latches_4_25(latches_4_25),
	.latches_4_26(latches_4_26),
	.latches_4_24(latches_4_24),
	.latches_5_15(latches_5_15),
	.latches_5_13(latches_5_13),
	.latches_5_14(latches_5_14),
	.latches_5_12(latches_5_12),
	.latches_5_11(latches_5_11),
	.latches_5_9(latches_5_9),
	.latches_5_10(latches_5_10),
	.latches_5_8(latches_5_8),
	.latches_5_1(latches_5_1),
	.latches_5_2(latches_5_2),
	.latches_5_0(latches_5_0),
	.latches_5_3(latches_5_3),
	.latches_5_21(latches_5_21),
	.latches_5_22(latches_5_22),
	.latches_5_20(latches_5_20),
	.latches_5_23(latches_5_23),
	.latches_5_17(latches_5_17),
	.latches_5_18(latches_5_18),
	.latches_5_16(latches_5_16),
	.latches_5_19(latches_5_19),
	.latches_5_5(latches_5_5),
	.latches_5_6(latches_5_6),
	.latches_5_4(latches_5_4),
	.latches_5_7(latches_5_7),
	.latches_5_31(latches_5_31),
	.latches_5_29(latches_5_29),
	.latches_5_30(latches_5_30),
	.latches_5_28(latches_5_28),
	.latches_5_27(latches_5_27),
	.latches_5_25(latches_5_25),
	.latches_5_26(latches_5_26),
	.latches_5_24(latches_5_24),
	.latches_6_15(latches_6_15),
	.latches_6_13(latches_6_13),
	.latches_6_14(latches_6_14),
	.latches_6_12(latches_6_12),
	.latches_6_11(latches_6_11),
	.latches_6_9(latches_6_9),
	.latches_6_10(latches_6_10),
	.latches_6_8(latches_6_8),
	.latches_6_1(latches_6_1),
	.latches_6_2(latches_6_2),
	.latches_6_0(latches_6_0),
	.latches_6_3(latches_6_3),
	.latches_6_21(latches_6_21),
	.latches_6_22(latches_6_22),
	.latches_6_20(latches_6_20),
	.latches_6_23(latches_6_23),
	.latches_6_17(latches_6_17),
	.latches_6_18(latches_6_18),
	.latches_6_16(latches_6_16),
	.latches_6_19(latches_6_19),
	.latches_6_5(latches_6_5),
	.latches_6_6(latches_6_6),
	.latches_6_4(latches_6_4),
	.latches_6_7(latches_6_7),
	.latches_6_31(latches_6_31),
	.latches_6_29(latches_6_29),
	.latches_6_30(latches_6_30),
	.latches_6_28(latches_6_28),
	.latches_6_27(latches_6_27),
	.latches_6_25(latches_6_25),
	.latches_6_26(latches_6_26),
	.latches_6_24(latches_6_24),
	.latches_7_15(latches_7_15),
	.latches_7_13(latches_7_13),
	.latches_7_14(latches_7_14),
	.latches_7_12(latches_7_12),
	.latches_7_11(latches_7_11),
	.latches_7_9(latches_7_9),
	.latches_7_10(latches_7_10),
	.latches_7_8(latches_7_8),
	.latches_7_1(latches_7_1),
	.latches_7_2(latches_7_2),
	.latches_7_0(latches_7_0),
	.latches_7_3(latches_7_3),
	.latches_7_21(latches_7_21),
	.latches_7_22(latches_7_22),
	.latches_7_20(latches_7_20),
	.latches_7_23(latches_7_23),
	.latches_7_17(latches_7_17),
	.latches_7_18(latches_7_18),
	.latches_7_16(latches_7_16),
	.latches_7_19(latches_7_19),
	.latches_7_5(latches_7_5),
	.latches_7_6(latches_7_6),
	.latches_7_4(latches_7_4),
	.latches_7_7(latches_7_7),
	.latches_7_31(latches_7_31),
	.latches_7_29(latches_7_29),
	.latches_7_30(latches_7_30),
	.latches_7_28(latches_7_28),
	.latches_7_27(latches_7_27),
	.latches_7_25(latches_7_25),
	.latches_7_26(latches_7_26),
	.latches_7_24(latches_7_24),
	.latches_8_15(latches_8_15),
	.latches_8_13(latches_8_13),
	.latches_8_14(latches_8_14),
	.latches_8_12(latches_8_12),
	.latches_8_11(latches_8_11),
	.latches_8_9(latches_8_9),
	.latches_8_10(latches_8_10),
	.latches_8_8(latches_8_8),
	.latches_8_1(latches_8_1),
	.latches_8_2(latches_8_2),
	.latches_8_0(latches_8_0),
	.latches_8_3(latches_8_3),
	.latches_8_21(latches_8_21),
	.latches_8_22(latches_8_22),
	.latches_8_20(latches_8_20),
	.latches_8_23(latches_8_23),
	.latches_8_17(latches_8_17),
	.latches_8_18(latches_8_18),
	.latches_8_16(latches_8_16),
	.latches_8_19(latches_8_19),
	.latches_8_5(latches_8_5),
	.latches_8_6(latches_8_6),
	.latches_8_4(latches_8_4),
	.latches_8_7(latches_8_7),
	.latches_8_31(latches_8_31),
	.latches_8_29(latches_8_29),
	.latches_8_30(latches_8_30),
	.latches_8_28(latches_8_28),
	.latches_8_27(latches_8_27),
	.latches_8_25(latches_8_25),
	.latches_8_26(latches_8_26),
	.latches_8_24(latches_8_24),
	.latches_9_15(latches_9_15),
	.latches_9_13(latches_9_13),
	.latches_9_14(latches_9_14),
	.latches_9_12(latches_9_12),
	.latches_9_11(latches_9_11),
	.latches_9_9(latches_9_9),
	.latches_9_10(latches_9_10),
	.latches_9_8(latches_9_8),
	.latches_9_1(latches_9_1),
	.latches_9_2(latches_9_2),
	.latches_9_0(latches_9_0),
	.latches_9_3(latches_9_3),
	.latches_9_21(latches_9_21),
	.latches_9_22(latches_9_22),
	.latches_9_20(latches_9_20),
	.latches_9_23(latches_9_23),
	.latches_9_17(latches_9_17),
	.latches_9_18(latches_9_18),
	.latches_9_16(latches_9_16),
	.latches_9_19(latches_9_19),
	.latches_9_5(latches_9_5),
	.latches_9_6(latches_9_6),
	.latches_9_4(latches_9_4),
	.latches_9_7(latches_9_7),
	.latches_9_31(latches_9_31),
	.latches_9_29(latches_9_29),
	.latches_9_30(latches_9_30),
	.latches_9_28(latches_9_28),
	.latches_9_27(latches_9_27),
	.latches_9_25(latches_9_25),
	.latches_9_26(latches_9_26),
	.latches_9_24(latches_9_24),
	.latches_10_15(latches_10_15),
	.latches_10_13(latches_10_13),
	.latches_10_14(latches_10_14),
	.latches_10_12(latches_10_12),
	.latches_10_11(latches_10_11),
	.latches_10_9(latches_10_9),
	.latches_10_10(latches_10_10),
	.latches_10_8(latches_10_8),
	.latches_10_1(latches_10_1),
	.latches_10_2(latches_10_2),
	.latches_10_0(latches_10_0),
	.latches_10_3(latches_10_3),
	.latches_10_21(latches_10_21),
	.latches_10_22(latches_10_22),
	.latches_10_20(latches_10_20),
	.latches_10_23(latches_10_23),
	.latches_10_17(latches_10_17),
	.latches_10_18(latches_10_18),
	.latches_10_16(latches_10_16),
	.latches_10_19(latches_10_19),
	.latches_10_5(latches_10_5),
	.latches_10_6(latches_10_6),
	.latches_10_4(latches_10_4),
	.latches_10_7(latches_10_7),
	.latches_10_31(latches_10_31),
	.latches_10_29(latches_10_29),
	.latches_10_30(latches_10_30),
	.latches_10_28(latches_10_28),
	.latches_10_27(latches_10_27),
	.latches_10_25(latches_10_25),
	.latches_10_26(latches_10_26),
	.latches_10_24(latches_10_24),
	.latches_11_15(latches_11_15),
	.latches_11_13(latches_11_13),
	.latches_11_14(latches_11_14),
	.latches_11_12(latches_11_12),
	.latches_11_11(latches_11_11),
	.latches_11_9(latches_11_9),
	.latches_11_10(latches_11_10),
	.latches_11_8(latches_11_8),
	.latches_11_1(latches_11_1),
	.latches_11_2(latches_11_2),
	.latches_11_0(latches_11_0),
	.latches_11_3(latches_11_3),
	.latches_11_21(latches_11_21),
	.latches_11_22(latches_11_22),
	.latches_11_20(latches_11_20),
	.latches_11_23(latches_11_23),
	.latches_11_17(latches_11_17),
	.latches_11_18(latches_11_18),
	.latches_11_16(latches_11_16),
	.latches_11_19(latches_11_19),
	.latches_11_5(latches_11_5),
	.latches_11_6(latches_11_6),
	.latches_11_4(latches_11_4),
	.latches_11_7(latches_11_7),
	.latches_11_31(latches_11_31),
	.latches_11_29(latches_11_29),
	.latches_11_30(latches_11_30),
	.latches_11_28(latches_11_28),
	.latches_11_27(latches_11_27),
	.latches_11_25(latches_11_25),
	.latches_11_26(latches_11_26),
	.latches_11_24(latches_11_24),
	.latches_12_15(latches_12_15),
	.latches_12_13(latches_12_13),
	.latches_12_14(latches_12_14),
	.latches_12_12(latches_12_12),
	.latches_12_11(latches_12_11),
	.latches_12_9(latches_12_9),
	.latches_12_10(latches_12_10),
	.latches_12_8(latches_12_8),
	.latches_12_1(latches_12_1),
	.latches_12_2(latches_12_2),
	.latches_12_0(latches_12_0),
	.latches_12_3(latches_12_3),
	.latches_12_21(latches_12_21),
	.latches_12_22(latches_12_22),
	.latches_12_20(latches_12_20),
	.latches_12_23(latches_12_23),
	.latches_12_17(latches_12_17),
	.latches_12_18(latches_12_18),
	.latches_12_16(latches_12_16),
	.latches_12_19(latches_12_19),
	.latches_12_5(latches_12_5),
	.latches_12_6(latches_12_6),
	.latches_12_4(latches_12_4),
	.latches_12_7(latches_12_7),
	.latches_12_31(latches_12_31),
	.latches_12_29(latches_12_29),
	.latches_12_30(latches_12_30),
	.latches_12_28(latches_12_28),
	.latches_12_27(latches_12_27),
	.latches_12_25(latches_12_25),
	.latches_12_26(latches_12_26),
	.latches_12_24(latches_12_24),
	.latches_13_15(latches_13_15),
	.latches_13_13(latches_13_13),
	.latches_13_14(latches_13_14),
	.latches_13_12(latches_13_12),
	.latches_13_11(latches_13_11),
	.latches_13_9(latches_13_9),
	.latches_13_10(latches_13_10),
	.latches_13_8(latches_13_8),
	.latches_13_1(latches_13_1),
	.latches_13_2(latches_13_2),
	.latches_13_0(latches_13_0),
	.latches_13_3(latches_13_3),
	.latches_13_21(latches_13_21),
	.latches_13_22(latches_13_22),
	.latches_13_20(latches_13_20),
	.latches_13_23(latches_13_23),
	.latches_13_17(latches_13_17),
	.latches_13_18(latches_13_18),
	.latches_13_16(latches_13_16),
	.latches_13_19(latches_13_19),
	.latches_13_5(latches_13_5),
	.latches_13_6(latches_13_6),
	.latches_13_4(latches_13_4),
	.latches_13_7(latches_13_7),
	.latches_13_31(latches_13_31),
	.latches_13_29(latches_13_29),
	.latches_13_30(latches_13_30),
	.latches_13_28(latches_13_28),
	.latches_13_27(latches_13_27),
	.latches_13_25(latches_13_25),
	.latches_13_26(latches_13_26),
	.latches_13_24(latches_13_24),
	.latches_14_15(latches_14_15),
	.latches_14_13(latches_14_13),
	.latches_14_14(latches_14_14),
	.latches_14_12(latches_14_12),
	.latches_14_11(latches_14_11),
	.latches_14_9(latches_14_9),
	.latches_14_10(latches_14_10),
	.latches_14_8(latches_14_8),
	.latches_14_1(latches_14_1),
	.latches_14_2(latches_14_2),
	.latches_14_0(latches_14_0),
	.latches_14_3(latches_14_3),
	.latches_14_21(latches_14_21),
	.latches_14_22(latches_14_22),
	.latches_14_20(latches_14_20),
	.latches_14_23(latches_14_23),
	.latches_14_17(latches_14_17),
	.latches_14_18(latches_14_18),
	.latches_14_16(latches_14_16),
	.latches_14_19(latches_14_19),
	.latches_14_5(latches_14_5),
	.latches_14_6(latches_14_6),
	.latches_14_4(latches_14_4),
	.latches_14_7(latches_14_7),
	.latches_14_31(latches_14_31),
	.latches_14_29(latches_14_29),
	.latches_14_30(latches_14_30),
	.latches_14_28(latches_14_28),
	.latches_14_27(latches_14_27),
	.latches_14_25(latches_14_25),
	.latches_14_26(latches_14_26),
	.latches_14_24(latches_14_24),
	.latches_15_15(latches_15_15),
	.latches_15_13(latches_15_13),
	.latches_15_14(latches_15_14),
	.latches_15_12(latches_15_12),
	.latches_15_11(latches_15_11),
	.latches_15_9(latches_15_9),
	.latches_15_10(latches_15_10),
	.latches_15_8(latches_15_8),
	.latches_15_1(latches_15_1),
	.latches_15_2(latches_15_2),
	.latches_15_0(latches_15_0),
	.latches_15_3(latches_15_3),
	.latches_15_21(latches_15_21),
	.latches_15_22(latches_15_22),
	.latches_15_20(latches_15_20),
	.latches_15_23(latches_15_23),
	.latches_15_17(latches_15_17),
	.latches_15_18(latches_15_18),
	.latches_15_16(latches_15_16),
	.latches_15_19(latches_15_19),
	.latches_15_5(latches_15_5),
	.latches_15_6(latches_15_6),
	.latches_15_4(latches_15_4),
	.latches_15_7(latches_15_7),
	.latches_15_31(latches_15_31),
	.latches_15_29(latches_15_29),
	.latches_15_30(latches_15_30),
	.latches_15_28(latches_15_28),
	.latches_15_27(latches_15_27),
	.latches_15_25(latches_15_25),
	.latches_15_26(latches_15_26),
	.latches_15_24(latches_15_24));

endmodule

module memory_mux_v9c (
	address_0,
	address_1,
	address_2,
	address_4,
	address_3,
	w_anode196w_2,
	w_anode287w_2,
	w_anode165w_3,
	w_anode155w_3,
	w_anode125w_3,
	w_anode114w_3,
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	latches_0_15,
	latches_0_13,
	latches_0_14,
	latches_0_12,
	latches_0_11,
	latches_0_9,
	latches_0_10,
	latches_0_8,
	latches_0_1,
	latches_0_2,
	latches_0_0,
	latches_0_3,
	latches_0_21,
	latches_0_22,
	latches_0_20,
	latches_0_23,
	latches_0_17,
	latches_0_18,
	latches_0_16,
	latches_0_19,
	latches_0_5,
	latches_0_6,
	latches_0_4,
	latches_0_7,
	latches_0_31,
	latches_0_29,
	latches_0_30,
	latches_0_28,
	latches_0_27,
	latches_0_25,
	latches_0_26,
	latches_0_24,
	latches_1_15,
	latches_1_13,
	latches_1_14,
	latches_1_12,
	latches_1_11,
	latches_1_9,
	latches_1_10,
	latches_1_8,
	latches_1_1,
	latches_1_2,
	latches_1_0,
	latches_1_3,
	latches_1_21,
	latches_1_22,
	latches_1_20,
	latches_1_23,
	latches_1_17,
	latches_1_18,
	latches_1_16,
	latches_1_19,
	latches_1_5,
	latches_1_6,
	latches_1_4,
	latches_1_7,
	latches_1_31,
	latches_1_29,
	latches_1_30,
	latches_1_28,
	latches_1_27,
	latches_1_25,
	latches_1_26,
	latches_1_24,
	latches_2_15,
	latches_2_13,
	latches_2_14,
	latches_2_12,
	latches_2_11,
	latches_2_9,
	latches_2_10,
	latches_2_8,
	latches_2_1,
	latches_2_2,
	latches_2_0,
	latches_2_3,
	latches_2_21,
	latches_2_22,
	latches_2_20,
	latches_2_23,
	latches_2_17,
	latches_2_18,
	latches_2_16,
	latches_2_19,
	latches_2_5,
	latches_2_6,
	latches_2_4,
	latches_2_7,
	latches_2_31,
	latches_2_29,
	latches_2_30,
	latches_2_28,
	latches_2_27,
	latches_2_25,
	latches_2_26,
	latches_2_24,
	latches_3_15,
	latches_3_13,
	latches_3_14,
	latches_3_12,
	latches_3_11,
	latches_3_9,
	latches_3_10,
	latches_3_8,
	latches_3_1,
	latches_3_2,
	latches_3_0,
	latches_3_3,
	latches_3_21,
	latches_3_22,
	latches_3_20,
	latches_3_23,
	latches_3_17,
	latches_3_18,
	latches_3_16,
	latches_3_19,
	latches_3_5,
	latches_3_6,
	latches_3_4,
	latches_3_7,
	latches_3_31,
	latches_3_29,
	latches_3_30,
	latches_3_28,
	latches_3_27,
	latches_3_25,
	latches_3_26,
	latches_3_24,
	latches_4_15,
	latches_4_13,
	latches_4_14,
	latches_4_12,
	latches_4_11,
	latches_4_9,
	latches_4_10,
	latches_4_8,
	latches_4_1,
	latches_4_2,
	latches_4_0,
	latches_4_3,
	latches_4_21,
	latches_4_22,
	latches_4_20,
	latches_4_23,
	latches_4_17,
	latches_4_18,
	latches_4_16,
	latches_4_19,
	latches_4_5,
	latches_4_6,
	latches_4_4,
	latches_4_7,
	latches_4_31,
	latches_4_29,
	latches_4_30,
	latches_4_28,
	latches_4_27,
	latches_4_25,
	latches_4_26,
	latches_4_24,
	latches_5_15,
	latches_5_13,
	latches_5_14,
	latches_5_12,
	latches_5_11,
	latches_5_9,
	latches_5_10,
	latches_5_8,
	latches_5_1,
	latches_5_2,
	latches_5_0,
	latches_5_3,
	latches_5_21,
	latches_5_22,
	latches_5_20,
	latches_5_23,
	latches_5_17,
	latches_5_18,
	latches_5_16,
	latches_5_19,
	latches_5_5,
	latches_5_6,
	latches_5_4,
	latches_5_7,
	latches_5_31,
	latches_5_29,
	latches_5_30,
	latches_5_28,
	latches_5_27,
	latches_5_25,
	latches_5_26,
	latches_5_24,
	latches_6_15,
	latches_6_13,
	latches_6_14,
	latches_6_12,
	latches_6_11,
	latches_6_9,
	latches_6_10,
	latches_6_8,
	latches_6_1,
	latches_6_2,
	latches_6_0,
	latches_6_3,
	latches_6_21,
	latches_6_22,
	latches_6_20,
	latches_6_23,
	latches_6_17,
	latches_6_18,
	latches_6_16,
	latches_6_19,
	latches_6_5,
	latches_6_6,
	latches_6_4,
	latches_6_7,
	latches_6_31,
	latches_6_29,
	latches_6_30,
	latches_6_28,
	latches_6_27,
	latches_6_25,
	latches_6_26,
	latches_6_24,
	latches_7_15,
	latches_7_13,
	latches_7_14,
	latches_7_12,
	latches_7_11,
	latches_7_9,
	latches_7_10,
	latches_7_8,
	latches_7_1,
	latches_7_2,
	latches_7_0,
	latches_7_3,
	latches_7_21,
	latches_7_22,
	latches_7_20,
	latches_7_23,
	latches_7_17,
	latches_7_18,
	latches_7_16,
	latches_7_19,
	latches_7_5,
	latches_7_6,
	latches_7_4,
	latches_7_7,
	latches_7_31,
	latches_7_29,
	latches_7_30,
	latches_7_28,
	latches_7_27,
	latches_7_25,
	latches_7_26,
	latches_7_24,
	latches_8_15,
	latches_8_13,
	latches_8_14,
	latches_8_12,
	latches_8_11,
	latches_8_9,
	latches_8_10,
	latches_8_8,
	latches_8_1,
	latches_8_2,
	latches_8_0,
	latches_8_3,
	latches_8_21,
	latches_8_22,
	latches_8_20,
	latches_8_23,
	latches_8_17,
	latches_8_18,
	latches_8_16,
	latches_8_19,
	latches_8_5,
	latches_8_6,
	latches_8_4,
	latches_8_7,
	latches_8_31,
	latches_8_29,
	latches_8_30,
	latches_8_28,
	latches_8_27,
	latches_8_25,
	latches_8_26,
	latches_8_24,
	latches_9_15,
	latches_9_13,
	latches_9_14,
	latches_9_12,
	latches_9_11,
	latches_9_9,
	latches_9_10,
	latches_9_8,
	latches_9_1,
	latches_9_2,
	latches_9_0,
	latches_9_3,
	latches_9_21,
	latches_9_22,
	latches_9_20,
	latches_9_23,
	latches_9_17,
	latches_9_18,
	latches_9_16,
	latches_9_19,
	latches_9_5,
	latches_9_6,
	latches_9_4,
	latches_9_7,
	latches_9_31,
	latches_9_29,
	latches_9_30,
	latches_9_28,
	latches_9_27,
	latches_9_25,
	latches_9_26,
	latches_9_24,
	latches_10_15,
	latches_10_13,
	latches_10_14,
	latches_10_12,
	latches_10_11,
	latches_10_9,
	latches_10_10,
	latches_10_8,
	latches_10_1,
	latches_10_2,
	latches_10_0,
	latches_10_3,
	latches_10_21,
	latches_10_22,
	latches_10_20,
	latches_10_23,
	latches_10_17,
	latches_10_18,
	latches_10_16,
	latches_10_19,
	latches_10_5,
	latches_10_6,
	latches_10_4,
	latches_10_7,
	latches_10_31,
	latches_10_29,
	latches_10_30,
	latches_10_28,
	latches_10_27,
	latches_10_25,
	latches_10_26,
	latches_10_24,
	latches_11_15,
	latches_11_13,
	latches_11_14,
	latches_11_12,
	latches_11_11,
	latches_11_9,
	latches_11_10,
	latches_11_8,
	latches_11_1,
	latches_11_2,
	latches_11_0,
	latches_11_3,
	latches_11_21,
	latches_11_22,
	latches_11_20,
	latches_11_23,
	latches_11_17,
	latches_11_18,
	latches_11_16,
	latches_11_19,
	latches_11_5,
	latches_11_6,
	latches_11_4,
	latches_11_7,
	latches_11_31,
	latches_11_29,
	latches_11_30,
	latches_11_28,
	latches_11_27,
	latches_11_25,
	latches_11_26,
	latches_11_24,
	latches_12_15,
	latches_12_13,
	latches_12_14,
	latches_12_12,
	latches_12_11,
	latches_12_9,
	latches_12_10,
	latches_12_8,
	latches_12_1,
	latches_12_2,
	latches_12_0,
	latches_12_3,
	latches_12_21,
	latches_12_22,
	latches_12_20,
	latches_12_23,
	latches_12_17,
	latches_12_18,
	latches_12_16,
	latches_12_19,
	latches_12_5,
	latches_12_6,
	latches_12_4,
	latches_12_7,
	latches_12_31,
	latches_12_29,
	latches_12_30,
	latches_12_28,
	latches_12_27,
	latches_12_25,
	latches_12_26,
	latches_12_24,
	latches_13_15,
	latches_13_13,
	latches_13_14,
	latches_13_12,
	latches_13_11,
	latches_13_9,
	latches_13_10,
	latches_13_8,
	latches_13_1,
	latches_13_2,
	latches_13_0,
	latches_13_3,
	latches_13_21,
	latches_13_22,
	latches_13_20,
	latches_13_23,
	latches_13_17,
	latches_13_18,
	latches_13_16,
	latches_13_19,
	latches_13_5,
	latches_13_6,
	latches_13_4,
	latches_13_7,
	latches_13_31,
	latches_13_29,
	latches_13_30,
	latches_13_28,
	latches_13_27,
	latches_13_25,
	latches_13_26,
	latches_13_24,
	latches_14_15,
	latches_14_13,
	latches_14_14,
	latches_14_12,
	latches_14_11,
	latches_14_9,
	latches_14_10,
	latches_14_8,
	latches_14_1,
	latches_14_2,
	latches_14_0,
	latches_14_3,
	latches_14_21,
	latches_14_22,
	latches_14_20,
	latches_14_23,
	latches_14_17,
	latches_14_18,
	latches_14_16,
	latches_14_19,
	latches_14_5,
	latches_14_6,
	latches_14_4,
	latches_14_7,
	latches_14_31,
	latches_14_29,
	latches_14_30,
	latches_14_28,
	latches_14_27,
	latches_14_25,
	latches_14_26,
	latches_14_24,
	latches_15_15,
	latches_15_13,
	latches_15_14,
	latches_15_12,
	latches_15_11,
	latches_15_9,
	latches_15_10,
	latches_15_8,
	latches_15_1,
	latches_15_2,
	latches_15_0,
	latches_15_3,
	latches_15_21,
	latches_15_22,
	latches_15_20,
	latches_15_23,
	latches_15_17,
	latches_15_18,
	latches_15_16,
	latches_15_19,
	latches_15_5,
	latches_15_6,
	latches_15_4,
	latches_15_7,
	latches_15_31,
	latches_15_29,
	latches_15_30,
	latches_15_28,
	latches_15_27,
	latches_15_25,
	latches_15_26,
	latches_15_24)/* synthesis synthesis_greybox=0 */;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_4;
input 	address_3;
input 	w_anode196w_2;
input 	w_anode287w_2;
input 	w_anode165w_3;
input 	w_anode155w_3;
input 	w_anode125w_3;
input 	w_anode114w_3;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
input 	latches_0_15;
input 	latches_0_13;
input 	latches_0_14;
input 	latches_0_12;
input 	latches_0_11;
input 	latches_0_9;
input 	latches_0_10;
input 	latches_0_8;
input 	latches_0_1;
input 	latches_0_2;
input 	latches_0_0;
input 	latches_0_3;
input 	latches_0_21;
input 	latches_0_22;
input 	latches_0_20;
input 	latches_0_23;
input 	latches_0_17;
input 	latches_0_18;
input 	latches_0_16;
input 	latches_0_19;
input 	latches_0_5;
input 	latches_0_6;
input 	latches_0_4;
input 	latches_0_7;
input 	latches_0_31;
input 	latches_0_29;
input 	latches_0_30;
input 	latches_0_28;
input 	latches_0_27;
input 	latches_0_25;
input 	latches_0_26;
input 	latches_0_24;
input 	latches_1_15;
input 	latches_1_13;
input 	latches_1_14;
input 	latches_1_12;
input 	latches_1_11;
input 	latches_1_9;
input 	latches_1_10;
input 	latches_1_8;
input 	latches_1_1;
input 	latches_1_2;
input 	latches_1_0;
input 	latches_1_3;
input 	latches_1_21;
input 	latches_1_22;
input 	latches_1_20;
input 	latches_1_23;
input 	latches_1_17;
input 	latches_1_18;
input 	latches_1_16;
input 	latches_1_19;
input 	latches_1_5;
input 	latches_1_6;
input 	latches_1_4;
input 	latches_1_7;
input 	latches_1_31;
input 	latches_1_29;
input 	latches_1_30;
input 	latches_1_28;
input 	latches_1_27;
input 	latches_1_25;
input 	latches_1_26;
input 	latches_1_24;
input 	latches_2_15;
input 	latches_2_13;
input 	latches_2_14;
input 	latches_2_12;
input 	latches_2_11;
input 	latches_2_9;
input 	latches_2_10;
input 	latches_2_8;
input 	latches_2_1;
input 	latches_2_2;
input 	latches_2_0;
input 	latches_2_3;
input 	latches_2_21;
input 	latches_2_22;
input 	latches_2_20;
input 	latches_2_23;
input 	latches_2_17;
input 	latches_2_18;
input 	latches_2_16;
input 	latches_2_19;
input 	latches_2_5;
input 	latches_2_6;
input 	latches_2_4;
input 	latches_2_7;
input 	latches_2_31;
input 	latches_2_29;
input 	latches_2_30;
input 	latches_2_28;
input 	latches_2_27;
input 	latches_2_25;
input 	latches_2_26;
input 	latches_2_24;
input 	latches_3_15;
input 	latches_3_13;
input 	latches_3_14;
input 	latches_3_12;
input 	latches_3_11;
input 	latches_3_9;
input 	latches_3_10;
input 	latches_3_8;
input 	latches_3_1;
input 	latches_3_2;
input 	latches_3_0;
input 	latches_3_3;
input 	latches_3_21;
input 	latches_3_22;
input 	latches_3_20;
input 	latches_3_23;
input 	latches_3_17;
input 	latches_3_18;
input 	latches_3_16;
input 	latches_3_19;
input 	latches_3_5;
input 	latches_3_6;
input 	latches_3_4;
input 	latches_3_7;
input 	latches_3_31;
input 	latches_3_29;
input 	latches_3_30;
input 	latches_3_28;
input 	latches_3_27;
input 	latches_3_25;
input 	latches_3_26;
input 	latches_3_24;
input 	latches_4_15;
input 	latches_4_13;
input 	latches_4_14;
input 	latches_4_12;
input 	latches_4_11;
input 	latches_4_9;
input 	latches_4_10;
input 	latches_4_8;
input 	latches_4_1;
input 	latches_4_2;
input 	latches_4_0;
input 	latches_4_3;
input 	latches_4_21;
input 	latches_4_22;
input 	latches_4_20;
input 	latches_4_23;
input 	latches_4_17;
input 	latches_4_18;
input 	latches_4_16;
input 	latches_4_19;
input 	latches_4_5;
input 	latches_4_6;
input 	latches_4_4;
input 	latches_4_7;
input 	latches_4_31;
input 	latches_4_29;
input 	latches_4_30;
input 	latches_4_28;
input 	latches_4_27;
input 	latches_4_25;
input 	latches_4_26;
input 	latches_4_24;
input 	latches_5_15;
input 	latches_5_13;
input 	latches_5_14;
input 	latches_5_12;
input 	latches_5_11;
input 	latches_5_9;
input 	latches_5_10;
input 	latches_5_8;
input 	latches_5_1;
input 	latches_5_2;
input 	latches_5_0;
input 	latches_5_3;
input 	latches_5_21;
input 	latches_5_22;
input 	latches_5_20;
input 	latches_5_23;
input 	latches_5_17;
input 	latches_5_18;
input 	latches_5_16;
input 	latches_5_19;
input 	latches_5_5;
input 	latches_5_6;
input 	latches_5_4;
input 	latches_5_7;
input 	latches_5_31;
input 	latches_5_29;
input 	latches_5_30;
input 	latches_5_28;
input 	latches_5_27;
input 	latches_5_25;
input 	latches_5_26;
input 	latches_5_24;
input 	latches_6_15;
input 	latches_6_13;
input 	latches_6_14;
input 	latches_6_12;
input 	latches_6_11;
input 	latches_6_9;
input 	latches_6_10;
input 	latches_6_8;
input 	latches_6_1;
input 	latches_6_2;
input 	latches_6_0;
input 	latches_6_3;
input 	latches_6_21;
input 	latches_6_22;
input 	latches_6_20;
input 	latches_6_23;
input 	latches_6_17;
input 	latches_6_18;
input 	latches_6_16;
input 	latches_6_19;
input 	latches_6_5;
input 	latches_6_6;
input 	latches_6_4;
input 	latches_6_7;
input 	latches_6_31;
input 	latches_6_29;
input 	latches_6_30;
input 	latches_6_28;
input 	latches_6_27;
input 	latches_6_25;
input 	latches_6_26;
input 	latches_6_24;
input 	latches_7_15;
input 	latches_7_13;
input 	latches_7_14;
input 	latches_7_12;
input 	latches_7_11;
input 	latches_7_9;
input 	latches_7_10;
input 	latches_7_8;
input 	latches_7_1;
input 	latches_7_2;
input 	latches_7_0;
input 	latches_7_3;
input 	latches_7_21;
input 	latches_7_22;
input 	latches_7_20;
input 	latches_7_23;
input 	latches_7_17;
input 	latches_7_18;
input 	latches_7_16;
input 	latches_7_19;
input 	latches_7_5;
input 	latches_7_6;
input 	latches_7_4;
input 	latches_7_7;
input 	latches_7_31;
input 	latches_7_29;
input 	latches_7_30;
input 	latches_7_28;
input 	latches_7_27;
input 	latches_7_25;
input 	latches_7_26;
input 	latches_7_24;
input 	latches_8_15;
input 	latches_8_13;
input 	latches_8_14;
input 	latches_8_12;
input 	latches_8_11;
input 	latches_8_9;
input 	latches_8_10;
input 	latches_8_8;
input 	latches_8_1;
input 	latches_8_2;
input 	latches_8_0;
input 	latches_8_3;
input 	latches_8_21;
input 	latches_8_22;
input 	latches_8_20;
input 	latches_8_23;
input 	latches_8_17;
input 	latches_8_18;
input 	latches_8_16;
input 	latches_8_19;
input 	latches_8_5;
input 	latches_8_6;
input 	latches_8_4;
input 	latches_8_7;
input 	latches_8_31;
input 	latches_8_29;
input 	latches_8_30;
input 	latches_8_28;
input 	latches_8_27;
input 	latches_8_25;
input 	latches_8_26;
input 	latches_8_24;
input 	latches_9_15;
input 	latches_9_13;
input 	latches_9_14;
input 	latches_9_12;
input 	latches_9_11;
input 	latches_9_9;
input 	latches_9_10;
input 	latches_9_8;
input 	latches_9_1;
input 	latches_9_2;
input 	latches_9_0;
input 	latches_9_3;
input 	latches_9_21;
input 	latches_9_22;
input 	latches_9_20;
input 	latches_9_23;
input 	latches_9_17;
input 	latches_9_18;
input 	latches_9_16;
input 	latches_9_19;
input 	latches_9_5;
input 	latches_9_6;
input 	latches_9_4;
input 	latches_9_7;
input 	latches_9_31;
input 	latches_9_29;
input 	latches_9_30;
input 	latches_9_28;
input 	latches_9_27;
input 	latches_9_25;
input 	latches_9_26;
input 	latches_9_24;
input 	latches_10_15;
input 	latches_10_13;
input 	latches_10_14;
input 	latches_10_12;
input 	latches_10_11;
input 	latches_10_9;
input 	latches_10_10;
input 	latches_10_8;
input 	latches_10_1;
input 	latches_10_2;
input 	latches_10_0;
input 	latches_10_3;
input 	latches_10_21;
input 	latches_10_22;
input 	latches_10_20;
input 	latches_10_23;
input 	latches_10_17;
input 	latches_10_18;
input 	latches_10_16;
input 	latches_10_19;
input 	latches_10_5;
input 	latches_10_6;
input 	latches_10_4;
input 	latches_10_7;
input 	latches_10_31;
input 	latches_10_29;
input 	latches_10_30;
input 	latches_10_28;
input 	latches_10_27;
input 	latches_10_25;
input 	latches_10_26;
input 	latches_10_24;
input 	latches_11_15;
input 	latches_11_13;
input 	latches_11_14;
input 	latches_11_12;
input 	latches_11_11;
input 	latches_11_9;
input 	latches_11_10;
input 	latches_11_8;
input 	latches_11_1;
input 	latches_11_2;
input 	latches_11_0;
input 	latches_11_3;
input 	latches_11_21;
input 	latches_11_22;
input 	latches_11_20;
input 	latches_11_23;
input 	latches_11_17;
input 	latches_11_18;
input 	latches_11_16;
input 	latches_11_19;
input 	latches_11_5;
input 	latches_11_6;
input 	latches_11_4;
input 	latches_11_7;
input 	latches_11_31;
input 	latches_11_29;
input 	latches_11_30;
input 	latches_11_28;
input 	latches_11_27;
input 	latches_11_25;
input 	latches_11_26;
input 	latches_11_24;
input 	latches_12_15;
input 	latches_12_13;
input 	latches_12_14;
input 	latches_12_12;
input 	latches_12_11;
input 	latches_12_9;
input 	latches_12_10;
input 	latches_12_8;
input 	latches_12_1;
input 	latches_12_2;
input 	latches_12_0;
input 	latches_12_3;
input 	latches_12_21;
input 	latches_12_22;
input 	latches_12_20;
input 	latches_12_23;
input 	latches_12_17;
input 	latches_12_18;
input 	latches_12_16;
input 	latches_12_19;
input 	latches_12_5;
input 	latches_12_6;
input 	latches_12_4;
input 	latches_12_7;
input 	latches_12_31;
input 	latches_12_29;
input 	latches_12_30;
input 	latches_12_28;
input 	latches_12_27;
input 	latches_12_25;
input 	latches_12_26;
input 	latches_12_24;
input 	latches_13_15;
input 	latches_13_13;
input 	latches_13_14;
input 	latches_13_12;
input 	latches_13_11;
input 	latches_13_9;
input 	latches_13_10;
input 	latches_13_8;
input 	latches_13_1;
input 	latches_13_2;
input 	latches_13_0;
input 	latches_13_3;
input 	latches_13_21;
input 	latches_13_22;
input 	latches_13_20;
input 	latches_13_23;
input 	latches_13_17;
input 	latches_13_18;
input 	latches_13_16;
input 	latches_13_19;
input 	latches_13_5;
input 	latches_13_6;
input 	latches_13_4;
input 	latches_13_7;
input 	latches_13_31;
input 	latches_13_29;
input 	latches_13_30;
input 	latches_13_28;
input 	latches_13_27;
input 	latches_13_25;
input 	latches_13_26;
input 	latches_13_24;
input 	latches_14_15;
input 	latches_14_13;
input 	latches_14_14;
input 	latches_14_12;
input 	latches_14_11;
input 	latches_14_9;
input 	latches_14_10;
input 	latches_14_8;
input 	latches_14_1;
input 	latches_14_2;
input 	latches_14_0;
input 	latches_14_3;
input 	latches_14_21;
input 	latches_14_22;
input 	latches_14_20;
input 	latches_14_23;
input 	latches_14_17;
input 	latches_14_18;
input 	latches_14_16;
input 	latches_14_19;
input 	latches_14_5;
input 	latches_14_6;
input 	latches_14_4;
input 	latches_14_7;
input 	latches_14_31;
input 	latches_14_29;
input 	latches_14_30;
input 	latches_14_28;
input 	latches_14_27;
input 	latches_14_25;
input 	latches_14_26;
input 	latches_14_24;
input 	latches_15_15;
input 	latches_15_13;
input 	latches_15_14;
input 	latches_15_12;
input 	latches_15_11;
input 	latches_15_9;
input 	latches_15_10;
input 	latches_15_8;
input 	latches_15_1;
input 	latches_15_2;
input 	latches_15_0;
input 	latches_15_3;
input 	latches_15_21;
input 	latches_15_22;
input 	latches_15_20;
input 	latches_15_23;
input 	latches_15_17;
input 	latches_15_18;
input 	latches_15_16;
input 	latches_15_19;
input 	latches_15_5;
input 	latches_15_6;
input 	latches_15_4;
input 	latches_15_7;
input 	latches_15_31;
input 	latches_15_29;
input 	latches_15_30;
input 	latches_15_28;
input 	latches_15_27;
input 	latches_15_25;
input 	latches_15_26;
input 	latches_15_24;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_ram_dq_component|sram|mux|auto_generated|_~0_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~1_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~2_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~3_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~4_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~5_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~6_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~7_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~8_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~9_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~10_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~11_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~12_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~13_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~14_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~15_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~16_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~17_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~18_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~19_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~20_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~21_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~22_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~23_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~24_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~25_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~26_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~27_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~28_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~29_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~30_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~31_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~32_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~33_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~34_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~35_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~36_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~37_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~38_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~39_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~40_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~41_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~42_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~43_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~44_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~45_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~46_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~47_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~48_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~49_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~50_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~51_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~52_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~53_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~54_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~55_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~56_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~57_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~58_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~59_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~60_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~61_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~62_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~63_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~64_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~65_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~66_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~67_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~68_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~69_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~70_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~71_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~72_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~73_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~74_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~75_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~76_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~77_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~78_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~79_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~80_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~81_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~82_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~83_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~84_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~85_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~86_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~87_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~88_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~89_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~90_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~91_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~92_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~93_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~94_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~95_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~96_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~97_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~98_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~99_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~100_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~101_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~102_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~103_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~104_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~105_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~106_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~107_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~108_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~109_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~110_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~111_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~112_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~113_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~114_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~115_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~116_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~117_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~118_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~119_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~120_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~121_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~122_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~123_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~124_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~125_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~126_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~127_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~128_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~129_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~130_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~131_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~132_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~133_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~134_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~135_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~136_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~137_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~138_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~139_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~140_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~141_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~142_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~143_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~144_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~145_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~146_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~147_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~148_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~149_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~150_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~151_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~152_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~153_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~154_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~155_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~156_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~157_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~158_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|_~159_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207_combout ;
wire \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208_combout ;


maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_0),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~14 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_1),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~27 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_2),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~40 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_3),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~53 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_4),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~66 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_5),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~79 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_6),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~92 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_7),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~105 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_8),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~118 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_9),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~131 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_10),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~144 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_11),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~157 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_12),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~170 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_13),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~183 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_14),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~196 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203_combout ),
	.datac(w_anode287w_2),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(result_node_15),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 .lut_mask = "feee";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~209 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~0 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_0_15),
	.datac(latches_0_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~0_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~0 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~0 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~0 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~0 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~0 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~0 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~1 (
	.clk(gnd),
	.dataa(latches_0_14),
	.datab(latches_0_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~1_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~1 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~1 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~1 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~1 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~1 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~1 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~0_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~1_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_0_11),
	.datac(latches_0_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 (
	.clk(gnd),
	.dataa(latches_0_10),
	.datab(latches_0_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~1_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~2_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~2 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_0_2),
	.datac(address_1),
	.datad(latches_0_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~2_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~2 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~2 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~2 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~2 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~2 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~2 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~3 (
	.clk(gnd),
	.dataa(latches_0_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~2_combout ),
	.datad(latches_0_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~3_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~3 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~3 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~3 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~3 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~3 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~3 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 (
	.clk(gnd),
	.dataa(vcc),
	.datab(vcc),
	.datac(address_2),
	.datad(address_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 .lut_mask = "000f";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~0_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~3_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~3_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~5 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~4 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_0_22),
	.datac(address_1),
	.datad(latches_0_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~4_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~4 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~4 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~4 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~4 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~4 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~4 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~5 (
	.clk(gnd),
	.dataa(latches_0_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~4_combout ),
	.datad(latches_0_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~5_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~5 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~5 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~5 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~5 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~5 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~5 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~6 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_0_18),
	.datac(address_1),
	.datad(latches_0_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~6_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~6 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~6 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~6 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~6 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~6 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~6 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~7 (
	.clk(gnd),
	.dataa(latches_0_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~6_combout ),
	.datad(latches_0_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~7_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~7 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~7 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~7 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~7 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~7 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~7 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~5_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~7_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~8 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_0_6),
	.datac(address_1),
	.datad(latches_0_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~8_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~8 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~8 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~8 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~8 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~8 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~8 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~9 (
	.clk(gnd),
	.dataa(latches_0_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~8_combout ),
	.datad(latches_0_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~9_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~9 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~9 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~9 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~9 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~9 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~9 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 (
	.clk(gnd),
	.dataa(address_2),
	.datab(vcc),
	.datac(address_3),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 .lut_mask = "000a";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~6_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~9_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~8 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_0_31),
	.datac(latches_0_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_0_30),
	.datac(latches_0_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_0_27),
	.datac(latches_0_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_0_26),
	.datac(latches_0_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~9_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~10_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~11_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~12_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~13 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~10 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_1_15),
	.datac(latches_1_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~10_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~10 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~10 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~10 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~10 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~10 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~10 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~11 (
	.clk(gnd),
	.dataa(latches_1_14),
	.datab(latches_1_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~11_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~11 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~11 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~11 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~11 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~11 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~11 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~10_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~11_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_1_11),
	.datac(latches_1_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 (
	.clk(gnd),
	.dataa(latches_1_10),
	.datab(latches_1_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~16_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~17_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~12 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_1_2),
	.datac(address_1),
	.datad(latches_1_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~12_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~12 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~12 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~12 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~12 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~12 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~12 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~13 (
	.clk(gnd),
	.dataa(latches_1_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~12_combout ),
	.datad(latches_1_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~13_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~13 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~13 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~13 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~13 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~13 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~13 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~15_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~18_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~13_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~19 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~14 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_1_22),
	.datac(address_1),
	.datad(latches_1_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~14_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~14 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~14 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~14 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~14 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~14 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~14 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~15 (
	.clk(gnd),
	.dataa(latches_1_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~14_combout ),
	.datad(latches_1_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~15_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~15 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~15 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~15 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~15 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~15 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~15 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~16 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_1_18),
	.datac(address_1),
	.datad(latches_1_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~16_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~16 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~16 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~16 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~16 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~16 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~16 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~17 (
	.clk(gnd),
	.dataa(latches_1_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~16_combout ),
	.datad(latches_1_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~17_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~17 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~17 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~17 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~17 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~17 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~17 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~15_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~17_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~18 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_1_6),
	.datac(address_1),
	.datad(latches_1_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~18_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~18 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~18 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~18 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~18 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~18 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~18 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~19 (
	.clk(gnd),
	.dataa(latches_1_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~18_combout ),
	.datad(latches_1_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~19_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~19 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~19 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~19 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~19 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~19 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~19 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~20_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~19_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~21 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_1_31),
	.datac(latches_1_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_1_30),
	.datac(latches_1_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_1_27),
	.datac(latches_1_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_1_26),
	.datac(latches_1_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~22_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~23_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~24_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~25_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[1]~26 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~20 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_2_15),
	.datac(latches_2_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~20_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~20 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~20 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~20 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~20 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~20 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~20 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~21 (
	.clk(gnd),
	.dataa(latches_2_14),
	.datab(latches_2_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~21_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~21 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~21 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~21 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~21 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~21 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~21 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~20_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~21_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_2_11),
	.datac(latches_2_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 (
	.clk(gnd),
	.dataa(latches_2_10),
	.datab(latches_2_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~29_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~30_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~22 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_2_2),
	.datac(address_1),
	.datad(latches_2_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~22_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~22 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~22 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~22 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~22 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~22 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~22 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~23 (
	.clk(gnd),
	.dataa(latches_2_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~22_combout ),
	.datad(latches_2_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~23_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~23 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~23 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~23 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~23 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~23 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~23 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~28_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~31_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~23_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~32 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~24 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_2_22),
	.datac(address_1),
	.datad(latches_2_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~24_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~24 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~24 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~24 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~24 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~24 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~24 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~25 (
	.clk(gnd),
	.dataa(latches_2_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~24_combout ),
	.datad(latches_2_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~25_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~25 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~25 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~25 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~25 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~25 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~25 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~26 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_2_18),
	.datac(address_1),
	.datad(latches_2_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~26_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~26 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~26 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~26 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~26 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~26 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~26 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~27 (
	.clk(gnd),
	.dataa(latches_2_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~26_combout ),
	.datad(latches_2_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~27_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~27 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~27 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~27 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~27 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~27 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~27 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~25_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~27_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~28 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_2_6),
	.datac(address_1),
	.datad(latches_2_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~28_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~28 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~28 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~28 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~28 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~28 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~28 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~29 (
	.clk(gnd),
	.dataa(latches_2_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~28_combout ),
	.datad(latches_2_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~29_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~29 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~29 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~29 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~29 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~29 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~29 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~33_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~29_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~34 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_2_31),
	.datac(latches_2_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_2_30),
	.datac(latches_2_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_2_27),
	.datac(latches_2_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_2_26),
	.datac(latches_2_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~35_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~36_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~37_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~38_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[2]~39 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~30 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_3_15),
	.datac(latches_3_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~30_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~30 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~30 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~30 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~30 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~30 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~30 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~31 (
	.clk(gnd),
	.dataa(latches_3_14),
	.datab(latches_3_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~31_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~31 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~31 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~31 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~31 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~31 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~31 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~30_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~31_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_3_11),
	.datac(latches_3_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 (
	.clk(gnd),
	.dataa(latches_3_10),
	.datab(latches_3_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~42_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~43_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~32 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_3_2),
	.datac(address_1),
	.datad(latches_3_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~32_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~32 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~32 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~32 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~32 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~32 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~32 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~33 (
	.clk(gnd),
	.dataa(latches_3_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~32_combout ),
	.datad(latches_3_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~33_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~33 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~33 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~33 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~33 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~33 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~33 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~41_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~44_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~33_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~45 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~34 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_3_22),
	.datac(address_1),
	.datad(latches_3_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~34_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~34 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~34 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~34 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~34 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~34 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~34 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~35 (
	.clk(gnd),
	.dataa(latches_3_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~34_combout ),
	.datad(latches_3_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~35_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~35 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~35 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~35 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~35 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~35 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~35 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~36 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_3_18),
	.datac(address_1),
	.datad(latches_3_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~36_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~36 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~36 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~36 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~36 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~36 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~36 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~37 (
	.clk(gnd),
	.dataa(latches_3_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~36_combout ),
	.datad(latches_3_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~37_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~37 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~37 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~37 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~37 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~37 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~37 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~35_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~37_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~38 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_3_6),
	.datac(address_1),
	.datad(latches_3_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~38_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~38 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~38 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~38 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~38 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~38 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~38 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~39 (
	.clk(gnd),
	.dataa(latches_3_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~38_combout ),
	.datad(latches_3_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~39_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~39 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~39 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~39 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~39 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~39 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~39 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~46_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~39_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~47 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_3_31),
	.datac(latches_3_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_3_30),
	.datac(latches_3_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_3_27),
	.datac(latches_3_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_3_26),
	.datac(latches_3_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~48_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~49_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~50_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~51_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[3]~52 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~40 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_4_15),
	.datac(latches_4_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~40_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~40 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~40 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~40 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~40 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~40 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~40 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~41 (
	.clk(gnd),
	.dataa(latches_4_14),
	.datab(latches_4_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~41_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~41 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~41 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~41 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~41 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~41 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~41 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~40_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~41_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_4_11),
	.datac(latches_4_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 (
	.clk(gnd),
	.dataa(latches_4_10),
	.datab(latches_4_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~55_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~56_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~42 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_4_2),
	.datac(address_1),
	.datad(latches_4_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~42_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~42 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~42 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~42 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~42 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~42 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~42 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~43 (
	.clk(gnd),
	.dataa(latches_4_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~42_combout ),
	.datad(latches_4_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~43_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~43 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~43 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~43 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~43 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~43 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~43 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~54_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~57_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~43_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~58 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~44 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_4_22),
	.datac(address_1),
	.datad(latches_4_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~44_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~44 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~44 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~44 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~44 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~44 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~44 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~45 (
	.clk(gnd),
	.dataa(latches_4_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~44_combout ),
	.datad(latches_4_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~45_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~45 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~45 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~45 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~45 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~45 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~45 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~46 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_4_18),
	.datac(address_1),
	.datad(latches_4_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~46_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~46 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~46 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~46 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~46 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~46 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~46 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~47 (
	.clk(gnd),
	.dataa(latches_4_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~46_combout ),
	.datad(latches_4_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~47_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~47 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~47 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~47 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~47 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~47 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~47 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~45_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~47_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~48 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_4_6),
	.datac(address_1),
	.datad(latches_4_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~48_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~48 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~48 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~48 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~48 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~48 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~48 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~49 (
	.clk(gnd),
	.dataa(latches_4_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~48_combout ),
	.datad(latches_4_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~49_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~49 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~49 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~49 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~49 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~49 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~49 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~59_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~49_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~60 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_4_31),
	.datac(latches_4_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_4_30),
	.datac(latches_4_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_4_27),
	.datac(latches_4_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_4_26),
	.datac(latches_4_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~61_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~62_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~63_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~64_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[4]~65 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~50 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_5_15),
	.datac(latches_5_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~50_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~50 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~50 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~50 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~50 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~50 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~50 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~51 (
	.clk(gnd),
	.dataa(latches_5_14),
	.datab(latches_5_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~51_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~51 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~51 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~51 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~51 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~51 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~51 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~50_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~51_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_5_11),
	.datac(latches_5_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 (
	.clk(gnd),
	.dataa(latches_5_10),
	.datab(latches_5_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~68_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~69_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~52 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_5_2),
	.datac(address_1),
	.datad(latches_5_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~52_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~52 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~52 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~52 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~52 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~52 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~52 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~53 (
	.clk(gnd),
	.dataa(latches_5_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~52_combout ),
	.datad(latches_5_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~53_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~53 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~53 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~53 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~53 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~53 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~53 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~67_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~70_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~53_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~71 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~54 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_5_22),
	.datac(address_1),
	.datad(latches_5_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~54_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~54 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~54 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~54 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~54 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~54 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~54 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~55 (
	.clk(gnd),
	.dataa(latches_5_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~54_combout ),
	.datad(latches_5_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~55_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~55 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~55 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~55 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~55 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~55 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~55 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~56 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_5_18),
	.datac(address_1),
	.datad(latches_5_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~56_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~56 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~56 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~56 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~56 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~56 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~56 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~57 (
	.clk(gnd),
	.dataa(latches_5_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~56_combout ),
	.datad(latches_5_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~57_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~57 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~57 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~57 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~57 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~57 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~57 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~55_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~57_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~58 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_5_6),
	.datac(address_1),
	.datad(latches_5_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~58_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~58 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~58 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~58 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~58 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~58 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~58 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~59 (
	.clk(gnd),
	.dataa(latches_5_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~58_combout ),
	.datad(latches_5_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~59_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~59 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~59 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~59 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~59 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~59 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~59 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~72_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~59_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~73 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_5_31),
	.datac(latches_5_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_5_30),
	.datac(latches_5_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_5_27),
	.datac(latches_5_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_5_26),
	.datac(latches_5_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~74_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~75_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~76_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~77_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[5]~78 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~60 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_6_15),
	.datac(latches_6_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~60_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~60 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~60 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~60 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~60 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~60 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~60 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~61 (
	.clk(gnd),
	.dataa(latches_6_14),
	.datab(latches_6_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~61_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~61 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~61 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~61 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~61 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~61 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~61 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~60_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~61_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_6_11),
	.datac(latches_6_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 (
	.clk(gnd),
	.dataa(latches_6_10),
	.datab(latches_6_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~81_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~82_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~62 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_6_2),
	.datac(address_1),
	.datad(latches_6_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~62_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~62 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~62 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~62 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~62 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~62 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~62 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~63 (
	.clk(gnd),
	.dataa(latches_6_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~62_combout ),
	.datad(latches_6_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~63_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~63 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~63 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~63 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~63 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~63 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~63 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~80_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~83_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~63_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~84 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~64 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_6_22),
	.datac(address_1),
	.datad(latches_6_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~64_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~64 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~64 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~64 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~64 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~64 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~64 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~65 (
	.clk(gnd),
	.dataa(latches_6_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~64_combout ),
	.datad(latches_6_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~65_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~65 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~65 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~65 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~65 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~65 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~65 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~66 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_6_18),
	.datac(address_1),
	.datad(latches_6_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~66_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~66 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~66 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~66 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~66 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~66 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~66 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~67 (
	.clk(gnd),
	.dataa(latches_6_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~66_combout ),
	.datad(latches_6_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~67_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~67 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~67 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~67 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~67 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~67 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~67 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~65_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~67_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~68 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_6_6),
	.datac(address_1),
	.datad(latches_6_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~68_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~68 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~68 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~68 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~68 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~68 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~68 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~69 (
	.clk(gnd),
	.dataa(latches_6_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~68_combout ),
	.datad(latches_6_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~69_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~69 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~69 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~69 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~69 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~69 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~69 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~85_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~69_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~86 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_6_31),
	.datac(latches_6_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_6_30),
	.datac(latches_6_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_6_27),
	.datac(latches_6_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_6_26),
	.datac(latches_6_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~87_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~88_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~89_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~90_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[6]~91 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~70 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_7_15),
	.datac(latches_7_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~70_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~70 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~70 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~70 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~70 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~70 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~70 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~71 (
	.clk(gnd),
	.dataa(latches_7_14),
	.datab(latches_7_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~71_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~71 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~71 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~71 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~71 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~71 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~71 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~70_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~71_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_7_11),
	.datac(latches_7_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 (
	.clk(gnd),
	.dataa(latches_7_10),
	.datab(latches_7_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~94_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~95_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~72 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_7_2),
	.datac(address_1),
	.datad(latches_7_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~72_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~72 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~72 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~72 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~72 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~72 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~72 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~73 (
	.clk(gnd),
	.dataa(latches_7_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~72_combout ),
	.datad(latches_7_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~73_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~73 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~73 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~73 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~73 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~73 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~73 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~93_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~96_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~73_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~97 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~74 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_7_22),
	.datac(address_1),
	.datad(latches_7_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~74_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~74 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~74 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~74 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~74 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~74 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~74 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~75 (
	.clk(gnd),
	.dataa(latches_7_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~74_combout ),
	.datad(latches_7_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~75_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~75 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~75 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~75 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~75 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~75 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~75 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~76 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_7_18),
	.datac(address_1),
	.datad(latches_7_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~76_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~76 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~76 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~76 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~76 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~76 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~76 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~77 (
	.clk(gnd),
	.dataa(latches_7_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~76_combout ),
	.datad(latches_7_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~77_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~77 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~77 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~77 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~77 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~77 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~77 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~75_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~77_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~78 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_7_6),
	.datac(address_1),
	.datad(latches_7_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~78_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~78 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~78 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~78 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~78 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~78 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~78 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~79 (
	.clk(gnd),
	.dataa(latches_7_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~78_combout ),
	.datad(latches_7_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~79_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~79 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~79 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~79 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~79 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~79 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~79 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~98_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~79_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~99 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_7_31),
	.datac(latches_7_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_7_30),
	.datac(latches_7_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_7_27),
	.datac(latches_7_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_7_26),
	.datac(latches_7_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~100_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~101_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~102_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~103_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[7]~104 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~80 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_8_15),
	.datac(latches_8_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~80_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~80 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~80 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~80 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~80 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~80 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~80 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~81 (
	.clk(gnd),
	.dataa(latches_8_14),
	.datab(latches_8_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~81_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~81 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~81 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~81 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~81 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~81 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~81 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~80_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~81_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_8_11),
	.datac(latches_8_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 (
	.clk(gnd),
	.dataa(latches_8_10),
	.datab(latches_8_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~107_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~108_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~82 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_8_2),
	.datac(address_1),
	.datad(latches_8_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~82_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~82 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~82 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~82 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~82 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~82 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~82 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~83 (
	.clk(gnd),
	.dataa(latches_8_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~82_combout ),
	.datad(latches_8_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~83_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~83 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~83 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~83 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~83 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~83 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~83 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~106_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~109_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~83_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~110 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~84 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_8_22),
	.datac(address_1),
	.datad(latches_8_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~84_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~84 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~84 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~84 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~84 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~84 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~84 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~85 (
	.clk(gnd),
	.dataa(latches_8_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~84_combout ),
	.datad(latches_8_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~85_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~85 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~85 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~85 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~85 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~85 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~85 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~86 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_8_18),
	.datac(address_1),
	.datad(latches_8_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~86_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~86 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~86 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~86 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~86 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~86 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~86 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~87 (
	.clk(gnd),
	.dataa(latches_8_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~86_combout ),
	.datad(latches_8_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~87_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~87 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~87 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~87 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~87 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~87 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~87 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~85_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~87_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~88 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_8_6),
	.datac(address_1),
	.datad(latches_8_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~88_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~88 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~88 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~88 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~88 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~88 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~88 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~89 (
	.clk(gnd),
	.dataa(latches_8_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~88_combout ),
	.datad(latches_8_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~89_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~89 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~89 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~89 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~89 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~89 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~89 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~111_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~89_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~112 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_8_31),
	.datac(latches_8_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_8_30),
	.datac(latches_8_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_8_27),
	.datac(latches_8_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_8_26),
	.datac(latches_8_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~113_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~114_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~115_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~116_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[8]~117 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~90 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_9_15),
	.datac(latches_9_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~90_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~90 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~90 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~90 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~90 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~90 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~90 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~91 (
	.clk(gnd),
	.dataa(latches_9_14),
	.datab(latches_9_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~91_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~91 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~91 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~91 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~91 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~91 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~91 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~90_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~91_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_9_11),
	.datac(latches_9_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 (
	.clk(gnd),
	.dataa(latches_9_10),
	.datab(latches_9_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~120_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~121_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~92 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_9_2),
	.datac(address_1),
	.datad(latches_9_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~92_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~92 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~92 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~92 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~92 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~92 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~92 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~93 (
	.clk(gnd),
	.dataa(latches_9_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~92_combout ),
	.datad(latches_9_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~93_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~93 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~93 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~93 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~93 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~93 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~93 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~119_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~122_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~93_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~123 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~94 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_9_22),
	.datac(address_1),
	.datad(latches_9_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~94_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~94 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~94 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~94 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~94 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~94 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~94 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~95 (
	.clk(gnd),
	.dataa(latches_9_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~94_combout ),
	.datad(latches_9_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~95_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~95 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~95 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~95 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~95 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~95 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~95 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~96 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_9_18),
	.datac(address_1),
	.datad(latches_9_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~96_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~96 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~96 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~96 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~96 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~96 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~96 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~97 (
	.clk(gnd),
	.dataa(latches_9_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~96_combout ),
	.datad(latches_9_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~97_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~97 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~97 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~97 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~97 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~97 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~97 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~95_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~97_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~98 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_9_6),
	.datac(address_1),
	.datad(latches_9_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~98_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~98 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~98 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~98 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~98 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~98 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~98 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~99 (
	.clk(gnd),
	.dataa(latches_9_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~98_combout ),
	.datad(latches_9_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~99_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~99 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~99 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~99 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~99 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~99 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~99 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~124_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~99_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~125 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_9_31),
	.datac(latches_9_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_9_30),
	.datac(latches_9_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_9_27),
	.datac(latches_9_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_9_26),
	.datac(latches_9_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~126_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~127_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~128_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~129_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[9]~130 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~100 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_10_15),
	.datac(latches_10_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~100_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~100 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~100 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~100 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~100 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~100 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~100 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~101 (
	.clk(gnd),
	.dataa(latches_10_14),
	.datab(latches_10_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~101_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~101 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~101 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~101 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~101 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~101 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~101 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~100_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~101_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_10_11),
	.datac(latches_10_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 (
	.clk(gnd),
	.dataa(latches_10_10),
	.datab(latches_10_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~133_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~134_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~102 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_10_2),
	.datac(address_1),
	.datad(latches_10_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~102_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~102 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~102 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~102 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~102 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~102 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~102 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~103 (
	.clk(gnd),
	.dataa(latches_10_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~102_combout ),
	.datad(latches_10_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~103_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~103 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~103 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~103 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~103 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~103 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~103 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~132_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~135_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~103_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~136 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~104 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_10_22),
	.datac(address_1),
	.datad(latches_10_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~104_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~104 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~104 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~104 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~104 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~104 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~104 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~105 (
	.clk(gnd),
	.dataa(latches_10_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~104_combout ),
	.datad(latches_10_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~105_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~105 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~105 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~105 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~105 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~105 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~105 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~106 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_10_18),
	.datac(address_1),
	.datad(latches_10_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~106_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~106 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~106 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~106 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~106 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~106 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~106 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~107 (
	.clk(gnd),
	.dataa(latches_10_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~106_combout ),
	.datad(latches_10_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~107_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~107 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~107 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~107 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~107 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~107 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~107 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~105_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~107_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~108 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_10_6),
	.datac(address_1),
	.datad(latches_10_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~108_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~108 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~108 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~108 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~108 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~108 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~108 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~109 (
	.clk(gnd),
	.dataa(latches_10_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~108_combout ),
	.datad(latches_10_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~109_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~109 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~109 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~109 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~109 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~109 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~109 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~137_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~109_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~138 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_10_31),
	.datac(latches_10_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_10_30),
	.datac(latches_10_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_10_27),
	.datac(latches_10_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_10_26),
	.datac(latches_10_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~139_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~140_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~141_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~142_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[10]~143 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~110 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_11_15),
	.datac(latches_11_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~110_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~110 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~110 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~110 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~110 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~110 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~110 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~111 (
	.clk(gnd),
	.dataa(latches_11_14),
	.datab(latches_11_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~111_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~111 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~111 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~111 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~111 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~111 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~111 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~110_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~111_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_11_11),
	.datac(latches_11_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 (
	.clk(gnd),
	.dataa(latches_11_10),
	.datab(latches_11_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~146_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~147_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~112 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_11_2),
	.datac(address_1),
	.datad(latches_11_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~112_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~112 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~112 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~112 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~112 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~112 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~112 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~113 (
	.clk(gnd),
	.dataa(latches_11_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~112_combout ),
	.datad(latches_11_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~113_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~113 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~113 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~113 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~113 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~113 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~113 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~145_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~148_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~113_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~149 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~114 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_11_22),
	.datac(address_1),
	.datad(latches_11_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~114_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~114 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~114 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~114 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~114 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~114 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~114 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~115 (
	.clk(gnd),
	.dataa(latches_11_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~114_combout ),
	.datad(latches_11_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~115_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~115 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~115 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~115 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~115 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~115 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~115 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~116 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_11_18),
	.datac(address_1),
	.datad(latches_11_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~116_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~116 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~116 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~116 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~116 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~116 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~116 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~117 (
	.clk(gnd),
	.dataa(latches_11_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~116_combout ),
	.datad(latches_11_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~117_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~117 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~117 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~117 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~117 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~117 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~117 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~115_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~117_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~118 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_11_6),
	.datac(address_1),
	.datad(latches_11_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~118_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~118 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~118 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~118 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~118 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~118 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~118 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~119 (
	.clk(gnd),
	.dataa(latches_11_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~118_combout ),
	.datad(latches_11_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~119_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~119 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~119 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~119 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~119 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~119 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~119 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~150_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~119_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~151 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_11_31),
	.datac(latches_11_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_11_30),
	.datac(latches_11_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_11_27),
	.datac(latches_11_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_11_26),
	.datac(latches_11_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~152_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~153_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~154_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~155_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[11]~156 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~120 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_12_15),
	.datac(latches_12_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~120_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~120 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~120 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~120 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~120 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~120 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~120 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~121 (
	.clk(gnd),
	.dataa(latches_12_14),
	.datab(latches_12_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~121_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~121 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~121 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~121 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~121 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~121 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~121 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~120_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~121_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_12_11),
	.datac(latches_12_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 (
	.clk(gnd),
	.dataa(latches_12_10),
	.datab(latches_12_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~159_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~160_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~122 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_12_2),
	.datac(address_1),
	.datad(latches_12_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~122_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~122 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~122 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~122 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~122 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~122 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~122 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~123 (
	.clk(gnd),
	.dataa(latches_12_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~122_combout ),
	.datad(latches_12_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~123_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~123 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~123 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~123 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~123 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~123 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~123 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~158_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~161_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~123_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~162 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~124 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_12_22),
	.datac(address_1),
	.datad(latches_12_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~124_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~124 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~124 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~124 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~124 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~124 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~124 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~125 (
	.clk(gnd),
	.dataa(latches_12_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~124_combout ),
	.datad(latches_12_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~125_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~125 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~125 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~125 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~125 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~125 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~125 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~126 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_12_18),
	.datac(address_1),
	.datad(latches_12_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~126_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~126 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~126 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~126 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~126 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~126 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~126 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~127 (
	.clk(gnd),
	.dataa(latches_12_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~126_combout ),
	.datad(latches_12_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~127_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~127 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~127 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~127 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~127 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~127 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~127 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~125_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~127_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~128 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_12_6),
	.datac(address_1),
	.datad(latches_12_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~128_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~128 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~128 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~128 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~128 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~128 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~128 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~129 (
	.clk(gnd),
	.dataa(latches_12_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~128_combout ),
	.datad(latches_12_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~129_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~129 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~129 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~129 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~129 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~129 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~129 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~163_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~129_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~164 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_12_31),
	.datac(latches_12_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_12_30),
	.datac(latches_12_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_12_27),
	.datac(latches_12_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_12_26),
	.datac(latches_12_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~165_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~166_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~167_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~168_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[12]~169 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~130 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_13_15),
	.datac(latches_13_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~130_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~130 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~130 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~130 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~130 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~130 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~130 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~131 (
	.clk(gnd),
	.dataa(latches_13_14),
	.datab(latches_13_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~131_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~131 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~131 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~131 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~131 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~131 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~131 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~130_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~131_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_13_11),
	.datac(latches_13_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 (
	.clk(gnd),
	.dataa(latches_13_10),
	.datab(latches_13_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~172_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~173_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~132 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_13_2),
	.datac(address_1),
	.datad(latches_13_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~132_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~132 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~132 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~132 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~132 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~132 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~132 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~133 (
	.clk(gnd),
	.dataa(latches_13_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~132_combout ),
	.datad(latches_13_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~133_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~133 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~133 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~133 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~133 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~133 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~133 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~171_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~174_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~133_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~175 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~134 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_13_22),
	.datac(address_1),
	.datad(latches_13_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~134_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~134 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~134 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~134 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~134 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~134 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~134 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~135 (
	.clk(gnd),
	.dataa(latches_13_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~134_combout ),
	.datad(latches_13_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~135_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~135 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~135 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~135 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~135 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~135 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~135 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~136 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_13_18),
	.datac(address_1),
	.datad(latches_13_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~136_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~136 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~136 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~136 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~136 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~136 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~136 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~137 (
	.clk(gnd),
	.dataa(latches_13_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~136_combout ),
	.datad(latches_13_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~137_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~137 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~137 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~137 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~137 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~137 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~137 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~135_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~137_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~138 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_13_6),
	.datac(address_1),
	.datad(latches_13_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~138_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~138 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~138 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~138 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~138 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~138 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~138 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~139 (
	.clk(gnd),
	.dataa(latches_13_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~138_combout ),
	.datad(latches_13_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~139_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~139 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~139 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~139 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~139 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~139 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~139 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~176_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~139_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~177 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_13_31),
	.datac(latches_13_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_13_30),
	.datac(latches_13_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_13_27),
	.datac(latches_13_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_13_26),
	.datac(latches_13_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~178_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~179_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~180_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~181_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[13]~182 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~140 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_14_15),
	.datac(latches_14_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~140_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~140 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~140 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~140 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~140 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~140 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~140 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~141 (
	.clk(gnd),
	.dataa(latches_14_14),
	.datab(latches_14_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~141_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~141 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~141 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~141 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~141 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~141 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~141 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~140_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~141_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_14_11),
	.datac(latches_14_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 (
	.clk(gnd),
	.dataa(latches_14_10),
	.datab(latches_14_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~185_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~186_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~142 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_14_2),
	.datac(address_1),
	.datad(latches_14_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~142_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~142 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~142 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~142 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~142 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~142 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~142 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~143 (
	.clk(gnd),
	.dataa(latches_14_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~142_combout ),
	.datad(latches_14_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~143_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~143 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~143 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~143 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~143 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~143 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~143 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~184_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~187_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~143_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~188 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~144 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_14_22),
	.datac(address_1),
	.datad(latches_14_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~144_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~144 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~144 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~144 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~144 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~144 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~144 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~145 (
	.clk(gnd),
	.dataa(latches_14_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~144_combout ),
	.datad(latches_14_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~145_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~145 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~145 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~145 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~145 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~145 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~145 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~146 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_14_18),
	.datac(address_1),
	.datad(latches_14_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~146_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~146 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~146 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~146 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~146 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~146 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~146 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~147 (
	.clk(gnd),
	.dataa(latches_14_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~146_combout ),
	.datad(latches_14_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~147_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~147 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~147 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~147 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~147 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~147 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~147 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~145_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~147_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~148 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_14_6),
	.datac(address_1),
	.datad(latches_14_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~148_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~148 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~148 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~148 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~148 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~148 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~148 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~149 (
	.clk(gnd),
	.dataa(latches_14_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~148_combout ),
	.datad(latches_14_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~149_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~149 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~149 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~149 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~149 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~149 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~149 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~189_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~149_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~190 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_14_31),
	.datac(latches_14_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_14_30),
	.datac(latches_14_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_14_27),
	.datac(latches_14_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_14_26),
	.datac(latches_14_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~191_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~192_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~193_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~194_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[14]~195 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~150 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_15_15),
	.datac(latches_15_13),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~150_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~150 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~150 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~150 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~150 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~150 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~150 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~151 (
	.clk(gnd),
	.dataa(latches_15_14),
	.datab(latches_15_12),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~151_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~151 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~151 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~151 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~151 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~151 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~151 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|_~150_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~151_combout ),
	.datac(address_2),
	.datad(address_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 .lut_mask = "00ef";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_15_11),
	.datac(latches_15_9),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 (
	.clk(gnd),
	.dataa(latches_15_10),
	.datab(latches_15_8),
	.datac(address_1),
	.datad(address_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 .lut_mask = "00ac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 (
	.clk(gnd),
	.dataa(address_3),
	.datab(address_2),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~198_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~199_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 .lut_mask = "aaa8";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~152 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_15_2),
	.datac(address_1),
	.datad(latches_15_0),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~152_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~152 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~152 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~152 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~152 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~152 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~152 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~153 (
	.clk(gnd),
	.dataa(latches_15_1),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~152_combout ),
	.datad(latches_15_3),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~153_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~153 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~153 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~153 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~153 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~153 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~153 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~197_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~200_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~4_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|_~153_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 .lut_mask = "a888";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~201 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~154 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_15_22),
	.datac(address_1),
	.datad(latches_15_20),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~154_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~154 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~154 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~154 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~154 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~154 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~154 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~155 (
	.clk(gnd),
	.dataa(latches_15_21),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~154_combout ),
	.datad(latches_15_23),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~155_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~155 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~155 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~155 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~155 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~155 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~155 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~156 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_15_18),
	.datac(address_1),
	.datad(latches_15_16),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~156_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~156 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~156 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~156 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~156 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~156 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~156 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~157 (
	.clk(gnd),
	.dataa(latches_15_17),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~156_combout ),
	.datad(latches_15_19),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~157_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~157 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~157 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~157 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~157 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~157 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~157 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 (
	.clk(gnd),
	.dataa(w_anode196w_2),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|_~155_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~157_combout ),
	.datad(address_2),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~158 (
	.clk(gnd),
	.dataa(address_0),
	.datab(latches_15_6),
	.datac(address_1),
	.datad(latches_15_4),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~158_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~158 .lut_mask = "e5e0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~158 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~158 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~158 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~158 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~158 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|_~159 (
	.clk(gnd),
	.dataa(latches_15_5),
	.datab(address_0),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~158_combout ),
	.datad(latches_15_7),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|_~159_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~159 .lut_mask = "f838";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~159 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~159 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~159 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~159 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|_~159 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~202_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[0]~7_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|_~159_combout ),
	.datad(vcc),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 .lut_mask = "eaea";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~203 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 (
	.clk(gnd),
	.dataa(w_anode165w_3),
	.datab(latches_15_31),
	.datac(latches_15_29),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 (
	.clk(gnd),
	.dataa(w_anode155w_3),
	.datab(latches_15_30),
	.datac(latches_15_28),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 (
	.clk(gnd),
	.dataa(w_anode125w_3),
	.datab(latches_15_27),
	.datac(latches_15_25),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 (
	.clk(gnd),
	.dataa(w_anode114w_3),
	.datab(latches_15_26),
	.datac(latches_15_24),
	.datad(address_1),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 .lut_mask = "88a0";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207 .synch_mode = "off";

maxv_lcell \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 (
	.clk(gnd),
	.dataa(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~204_combout ),
	.datab(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~205_combout ),
	.datac(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~206_combout ),
	.datad(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~207_combout ),
	.aclr(gnd),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.cin(gnd),
	.cin0(gnd),
	.cin1(vcc),
	.inverta(gnd),
	.regcascin(gnd),
	.combout(\lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208_combout ),
	.regout(),
	.cout(),
	.cout0(),
	.cout1());
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 .lut_mask = "fffe";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 .operation_mode = "normal";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 .output_mode = "comb_only";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 .register_cascade_mode = "off";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 .sum_lutc_input = "datac";
defparam \lpm_ram_dq_component|sram|mux|auto_generated|result_node[15]~208 .synch_mode = "off";

endmodule
